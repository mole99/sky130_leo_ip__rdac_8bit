** sch_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__rdac_8bit/xschem/sky130_leo_ip__rdac_8bit.sch
.subckt sky130_leo_ip__rdac_8bit D0 OUT D1 D2 D3 D4 D5 D6 D7 VGND
*.PININFO VGND:B D7:I D6:I D5:I D4:I D3:I D2:I D1:I D0:I OUT:O
XR1 D7 net1 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR2 net1 OUT VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR3 OUT net2 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR4 D6 net3 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR5 net3 net2 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR6 net2 net4 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR7 D5 net5 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR8 net5 net4 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR9 net4 net6 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR10 D4 net7 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR11 net7 net6 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR12 net6 net8 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR13 D3 net9 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR14 net9 net8 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR15 net8 net10 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR16 D2 net11 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR17 net11 net10 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR18 net10 net12 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR19 D1 net13 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR20 net13 net12 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR21 net12 net14 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR22 D0 net15 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR23 net15 net14 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR24 net14 net16 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR25 net16 VGND VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR26 VGND VGND VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR27 VGND VGND VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
**** begin user architecture code


* https://skywater-pdk.readthedocs.io/en/main/rules/device-details.html#p-poly-precision-resistors


**** end user architecture code
.ends
.end
