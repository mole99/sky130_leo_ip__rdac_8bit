* NGSPICE file created from sky130_leo_ip__rdac_8bit.ext - technology: sky130A

.subckt sky130_leo_ip__rdac_8bit D0 OUT D1 D2 D3 D4 D5 D6 D7 VGND
X0 a_6632_10921# a_6994_493# VGND.t30 sky130_fd_pr__res_high_po_1p41 l=50.12
X1 a_2288_10921# a_1202_10921# VGND.t20 sky130_fd_pr__res_high_po_1p41 l=50.12
X2 a_3374_10921# a_2288_10921# VGND.t28 sky130_fd_pr__res_high_po_1p41 l=50.12
X3 a_4460_10921# a_3374_10921# VGND.t29 sky130_fd_pr__res_high_po_1p41 l=50.12
X4 a_5546_10921# a_4460_10921# VGND.t22 sky130_fd_pr__res_high_po_1p41 l=50.12
X5 a_6632_10921# a_5546_10921# VGND.t13 sky130_fd_pr__res_high_po_1p41 l=50.12
X6 D1.t0 a_2650_493# VGND.t19 sky130_fd_pr__res_high_po_1p41 l=50.12
X7 a_7718_10921# a_6632_10921# VGND.t4 sky130_fd_pr__res_high_po_1p41 l=50.12
X8 OUT.t0 a_7718_10921# VGND.t0 sky130_fd_pr__res_high_po_1p41 l=50.12
X9 a_1202_10921# a_1564_493# VGND.t12 sky130_fd_pr__res_high_po_1p41 l=50.12
X10 a_2288_10921# a_2650_493# VGND.t11 sky130_fd_pr__res_high_po_1p41 l=50.12
X11 a_3374_10921# a_3736_493# VGND.t7 sky130_fd_pr__res_high_po_1p41 l=50.12
X12 a_4460_10921# a_4822_493# VGND.t27 sky130_fd_pr__res_high_po_1p41 l=50.12
X13 a_1202_10921# a_840_493# VGND.t31 sky130_fd_pr__res_high_po_1p41 l=50.12
X14 a_5546_10921# a_5908_493# VGND.t1 sky130_fd_pr__res_high_po_1p41 l=50.12
X15 VGND.t18 a_1564_493# VGND.t17 sky130_fd_pr__res_high_po_1p41 l=50.12
X16 a_7718_10921# a_8080_493# VGND.t2 sky130_fd_pr__res_high_po_1p41 l=50.12
X17 OUT.t1 a_9166_493# VGND.t6 sky130_fd_pr__res_high_po_1p41 l=50.12
X18 VGND.t24 VGND.t25 VGND.t23 sky130_fd_pr__res_high_po_1p41 l=50.12
X19 VGND.t9 VGND.t10 VGND.t8 sky130_fd_pr__res_high_po_1p41 l=50.12
X20 D2.t0 a_3736_493# VGND.t16 sky130_fd_pr__res_high_po_1p41 l=50.12
X21 D3.t0 a_4822_493# VGND.t15 sky130_fd_pr__res_high_po_1p41 l=50.12
X22 D4.t0 a_5908_493# VGND.t26 sky130_fd_pr__res_high_po_1p41 l=50.12
X23 D5.t0 a_6994_493# VGND.t3 sky130_fd_pr__res_high_po_1p41 l=50.12
X24 D6.t0 a_8080_493# VGND.t14 sky130_fd_pr__res_high_po_1p41 l=50.12
X25 D0.t0 a_840_493# VGND.t5 sky130_fd_pr__res_high_po_1p41 l=50.12
X26 D7.t0 a_9166_493# VGND.t21 sky130_fd_pr__res_high_po_1p41 l=50.12
R0 VGND.n1098 VGND.n626 585
R1 VGND.n1098 VGND.n632 585
R2 VGND.n1099 VGND.n1098 585
R3 VGND.n633 VGND.n632 585
R4 VGND.n1099 VGND.n633 585
R5 VGND.n860 VGND.n632 585
R6 VGND.n1099 VGND.n860 585
R7 VGND.n634 VGND.n632 585
R8 VGND.n1099 VGND.n634 585
R9 VGND.n858 VGND.n632 585
R10 VGND.n1099 VGND.n858 585
R11 VGND.n635 VGND.n632 585
R12 VGND.n1099 VGND.n635 585
R13 VGND.n856 VGND.n632 585
R14 VGND.n1099 VGND.n856 585
R15 VGND.n636 VGND.n632 585
R16 VGND.n1099 VGND.n636 585
R17 VGND.n854 VGND.n632 585
R18 VGND.n1099 VGND.n854 585
R19 VGND.n637 VGND.n632 585
R20 VGND.n1099 VGND.n637 585
R21 VGND.n852 VGND.n632 585
R22 VGND.n1099 VGND.n852 585
R23 VGND.n638 VGND.n632 585
R24 VGND.n1099 VGND.n638 585
R25 VGND.n850 VGND.n632 585
R26 VGND.n1099 VGND.n850 585
R27 VGND.n639 VGND.n632 585
R28 VGND.n1099 VGND.n639 585
R29 VGND.n848 VGND.n632 585
R30 VGND.n1099 VGND.n848 585
R31 VGND.n640 VGND.n632 585
R32 VGND.n1099 VGND.n640 585
R33 VGND.n846 VGND.n632 585
R34 VGND.n1099 VGND.n846 585
R35 VGND.n641 VGND.n632 585
R36 VGND.n1099 VGND.n641 585
R37 VGND.n844 VGND.n632 585
R38 VGND.n1099 VGND.n844 585
R39 VGND.n642 VGND.n632 585
R40 VGND.n1099 VGND.n642 585
R41 VGND.n842 VGND.n632 585
R42 VGND.n1099 VGND.n842 585
R43 VGND.n643 VGND.n632 585
R44 VGND.n1099 VGND.n643 585
R45 VGND.n840 VGND.n632 585
R46 VGND.n1099 VGND.n840 585
R47 VGND.n644 VGND.n632 585
R48 VGND.n1099 VGND.n644 585
R49 VGND.n838 VGND.n632 585
R50 VGND.n1099 VGND.n838 585
R51 VGND.n645 VGND.n632 585
R52 VGND.n1099 VGND.n645 585
R53 VGND.n836 VGND.n632 585
R54 VGND.n1099 VGND.n836 585
R55 VGND.n646 VGND.n632 585
R56 VGND.n1099 VGND.n646 585
R57 VGND.n834 VGND.n632 585
R58 VGND.n1099 VGND.n834 585
R59 VGND.n647 VGND.n632 585
R60 VGND.n1099 VGND.n647 585
R61 VGND.n832 VGND.n632 585
R62 VGND.n1099 VGND.n832 585
R63 VGND.n648 VGND.n632 585
R64 VGND.n1099 VGND.n648 585
R65 VGND.n830 VGND.n632 585
R66 VGND.n1099 VGND.n830 585
R67 VGND.n649 VGND.n632 585
R68 VGND.n1099 VGND.n649 585
R69 VGND.n828 VGND.n632 585
R70 VGND.n1099 VGND.n828 585
R71 VGND.n650 VGND.n632 585
R72 VGND.n1099 VGND.n650 585
R73 VGND.n826 VGND.n632 585
R74 VGND.n1099 VGND.n826 585
R75 VGND.n651 VGND.n632 585
R76 VGND.n1099 VGND.n651 585
R77 VGND.n824 VGND.n632 585
R78 VGND.n1099 VGND.n824 585
R79 VGND.n652 VGND.n632 585
R80 VGND.n1099 VGND.n652 585
R81 VGND.n822 VGND.n632 585
R82 VGND.n1099 VGND.n822 585
R83 VGND.n653 VGND.n632 585
R84 VGND.n1099 VGND.n653 585
R85 VGND.n820 VGND.n632 585
R86 VGND.n1099 VGND.n820 585
R87 VGND.n654 VGND.n632 585
R88 VGND.n1099 VGND.n654 585
R89 VGND.n818 VGND.n632 585
R90 VGND.n1099 VGND.n818 585
R91 VGND.n655 VGND.n632 585
R92 VGND.n1099 VGND.n655 585
R93 VGND.n816 VGND.n632 585
R94 VGND.n1099 VGND.n816 585
R95 VGND.n656 VGND.n632 585
R96 VGND.n1099 VGND.n656 585
R97 VGND.n814 VGND.n632 585
R98 VGND.n1099 VGND.n814 585
R99 VGND.n657 VGND.n632 585
R100 VGND.n1099 VGND.n657 585
R101 VGND.n812 VGND.n632 585
R102 VGND.n1099 VGND.n812 585
R103 VGND.n658 VGND.n632 585
R104 VGND.n1099 VGND.n658 585
R105 VGND.n810 VGND.n632 585
R106 VGND.n1099 VGND.n810 585
R107 VGND.n659 VGND.n632 585
R108 VGND.n1099 VGND.n659 585
R109 VGND.n808 VGND.n632 585
R110 VGND.n1099 VGND.n808 585
R111 VGND.n660 VGND.n632 585
R112 VGND.n1099 VGND.n660 585
R113 VGND.n806 VGND.n632 585
R114 VGND.n1099 VGND.n806 585
R115 VGND.n661 VGND.n632 585
R116 VGND.n1099 VGND.n661 585
R117 VGND.n804 VGND.n632 585
R118 VGND.n1099 VGND.n804 585
R119 VGND.n662 VGND.n632 585
R120 VGND.n1099 VGND.n662 585
R121 VGND.n802 VGND.n632 585
R122 VGND.n1099 VGND.n802 585
R123 VGND.n663 VGND.n632 585
R124 VGND.n1099 VGND.n663 585
R125 VGND.n800 VGND.n632 585
R126 VGND.n1099 VGND.n800 585
R127 VGND.n664 VGND.n632 585
R128 VGND.n1099 VGND.n664 585
R129 VGND.n798 VGND.n632 585
R130 VGND.n1099 VGND.n798 585
R131 VGND.n665 VGND.n632 585
R132 VGND.n1099 VGND.n665 585
R133 VGND.n796 VGND.n632 585
R134 VGND.n1099 VGND.n796 585
R135 VGND.n666 VGND.n632 585
R136 VGND.n1099 VGND.n666 585
R137 VGND.n794 VGND.n632 585
R138 VGND.n1099 VGND.n794 585
R139 VGND.n667 VGND.n632 585
R140 VGND.n1099 VGND.n667 585
R141 VGND.n792 VGND.n632 585
R142 VGND.n1099 VGND.n792 585
R143 VGND.n668 VGND.n632 585
R144 VGND.n1099 VGND.n668 585
R145 VGND.n790 VGND.n632 585
R146 VGND.n1099 VGND.n790 585
R147 VGND.n669 VGND.n632 585
R148 VGND.n1099 VGND.n669 585
R149 VGND.n788 VGND.n632 585
R150 VGND.n1099 VGND.n788 585
R151 VGND.n670 VGND.n632 585
R152 VGND.n1099 VGND.n670 585
R153 VGND.n786 VGND.n632 585
R154 VGND.n1099 VGND.n786 585
R155 VGND.n671 VGND.n632 585
R156 VGND.n1099 VGND.n671 585
R157 VGND.n784 VGND.n632 585
R158 VGND.n1099 VGND.n784 585
R159 VGND.n672 VGND.n632 585
R160 VGND.n1099 VGND.n672 585
R161 VGND.n782 VGND.n632 585
R162 VGND.n1099 VGND.n782 585
R163 VGND.n673 VGND.n632 585
R164 VGND.n1099 VGND.n673 585
R165 VGND.n780 VGND.n632 585
R166 VGND.n1099 VGND.n780 585
R167 VGND.n674 VGND.n632 585
R168 VGND.n1099 VGND.n674 585
R169 VGND.n778 VGND.n632 585
R170 VGND.n1099 VGND.n778 585
R171 VGND.n675 VGND.n632 585
R172 VGND.n1099 VGND.n675 585
R173 VGND.n776 VGND.n632 585
R174 VGND.n1099 VGND.n776 585
R175 VGND.n676 VGND.n632 585
R176 VGND.n1099 VGND.n676 585
R177 VGND.n774 VGND.n632 585
R178 VGND.n1099 VGND.n774 585
R179 VGND.n677 VGND.n632 585
R180 VGND.n1099 VGND.n677 585
R181 VGND.n772 VGND.n632 585
R182 VGND.n1099 VGND.n772 585
R183 VGND.n678 VGND.n632 585
R184 VGND.n1099 VGND.n678 585
R185 VGND.n770 VGND.n632 585
R186 VGND.n1099 VGND.n770 585
R187 VGND.n679 VGND.n632 585
R188 VGND.n1099 VGND.n679 585
R189 VGND.n768 VGND.n632 585
R190 VGND.n1099 VGND.n768 585
R191 VGND.n680 VGND.n632 585
R192 VGND.n1099 VGND.n680 585
R193 VGND.n766 VGND.n632 585
R194 VGND.n1099 VGND.n766 585
R195 VGND.n681 VGND.n632 585
R196 VGND.n1099 VGND.n681 585
R197 VGND.n764 VGND.n632 585
R198 VGND.n1099 VGND.n764 585
R199 VGND.n682 VGND.n632 585
R200 VGND.n1099 VGND.n682 585
R201 VGND.n762 VGND.n632 585
R202 VGND.n1099 VGND.n762 585
R203 VGND.n683 VGND.n632 585
R204 VGND.n1099 VGND.n683 585
R205 VGND.n760 VGND.n632 585
R206 VGND.n1099 VGND.n760 585
R207 VGND.n684 VGND.n632 585
R208 VGND.n1099 VGND.n684 585
R209 VGND.n758 VGND.n632 585
R210 VGND.n1099 VGND.n758 585
R211 VGND.n685 VGND.n632 585
R212 VGND.n1099 VGND.n685 585
R213 VGND.n756 VGND.n632 585
R214 VGND.n1099 VGND.n756 585
R215 VGND.n686 VGND.n632 585
R216 VGND.n1099 VGND.n686 585
R217 VGND.n754 VGND.n632 585
R218 VGND.n1099 VGND.n754 585
R219 VGND.n687 VGND.n632 585
R220 VGND.n1099 VGND.n687 585
R221 VGND.n752 VGND.n632 585
R222 VGND.n1099 VGND.n752 585
R223 VGND.n688 VGND.n632 585
R224 VGND.n1099 VGND.n688 585
R225 VGND.n750 VGND.n632 585
R226 VGND.n1099 VGND.n750 585
R227 VGND.n689 VGND.n632 585
R228 VGND.n1099 VGND.n689 585
R229 VGND.n748 VGND.n632 585
R230 VGND.n1099 VGND.n748 585
R231 VGND.n690 VGND.n632 585
R232 VGND.n1099 VGND.n690 585
R233 VGND.n746 VGND.n632 585
R234 VGND.n1099 VGND.n746 585
R235 VGND.n691 VGND.n632 585
R236 VGND.n1099 VGND.n691 585
R237 VGND.n744 VGND.n632 585
R238 VGND.n1099 VGND.n744 585
R239 VGND.n692 VGND.n632 585
R240 VGND.n1099 VGND.n692 585
R241 VGND.n742 VGND.n632 585
R242 VGND.n1099 VGND.n742 585
R243 VGND.n693 VGND.n632 585
R244 VGND.n1099 VGND.n693 585
R245 VGND.n740 VGND.n632 585
R246 VGND.n1099 VGND.n740 585
R247 VGND.n694 VGND.n632 585
R248 VGND.n1099 VGND.n694 585
R249 VGND.n738 VGND.n632 585
R250 VGND.n1099 VGND.n738 585
R251 VGND.n695 VGND.n632 585
R252 VGND.n1099 VGND.n695 585
R253 VGND.n736 VGND.n632 585
R254 VGND.n1099 VGND.n736 585
R255 VGND.n696 VGND.n632 585
R256 VGND.n1099 VGND.n696 585
R257 VGND.n734 VGND.n632 585
R258 VGND.n1099 VGND.n734 585
R259 VGND.n697 VGND.n632 585
R260 VGND.n1099 VGND.n697 585
R261 VGND.n732 VGND.n632 585
R262 VGND.n1099 VGND.n732 585
R263 VGND.n698 VGND.n632 585
R264 VGND.n1099 VGND.n698 585
R265 VGND.n730 VGND.n632 585
R266 VGND.n1099 VGND.n730 585
R267 VGND.n699 VGND.n632 585
R268 VGND.n1099 VGND.n699 585
R269 VGND.n728 VGND.n632 585
R270 VGND.n1099 VGND.n728 585
R271 VGND.n700 VGND.n632 585
R272 VGND.n1099 VGND.n700 585
R273 VGND.n726 VGND.n632 585
R274 VGND.n1099 VGND.n726 585
R275 VGND.n701 VGND.n632 585
R276 VGND.n1099 VGND.n701 585
R277 VGND.n724 VGND.n632 585
R278 VGND.n1099 VGND.n724 585
R279 VGND.n702 VGND.n632 585
R280 VGND.n1099 VGND.n702 585
R281 VGND.n722 VGND.n632 585
R282 VGND.n1099 VGND.n722 585
R283 VGND.n703 VGND.n632 585
R284 VGND.n1099 VGND.n703 585
R285 VGND.n720 VGND.n632 585
R286 VGND.n1099 VGND.n720 585
R287 VGND.n704 VGND.n632 585
R288 VGND.n1099 VGND.n704 585
R289 VGND.n718 VGND.n632 585
R290 VGND.n1099 VGND.n718 585
R291 VGND.n705 VGND.n632 585
R292 VGND.n1099 VGND.n705 585
R293 VGND.n716 VGND.n632 585
R294 VGND.n1099 VGND.n716 585
R295 VGND.n706 VGND.n632 585
R296 VGND.n1099 VGND.n706 585
R297 VGND.n714 VGND.n632 585
R298 VGND.n1099 VGND.n714 585
R299 VGND.n707 VGND.n632 585
R300 VGND.n1099 VGND.n707 585
R301 VGND.n712 VGND.n632 585
R302 VGND.n1099 VGND.n712 585
R303 VGND.n708 VGND.n632 585
R304 VGND.n1099 VGND.n708 585
R305 VGND.n710 VGND.n632 585
R306 VGND.n1099 VGND.n710 585
R307 VGND.n1100 VGND.n626 585
R308 VGND.n1100 VGND.n632 585
R309 VGND.n1100 VGND.n1099 585
R310 VGND.n180 VGND.n103 585
R311 VGND.n1561 VGND.n180 585
R312 VGND.n180 VGND.n97 585
R313 VGND.n1561 VGND.n184 585
R314 VGND.n184 VGND.n97 585
R315 VGND.n1561 VGND.n179 585
R316 VGND.n179 VGND.n97 585
R317 VGND.n1561 VGND.n187 585
R318 VGND.n187 VGND.n97 585
R319 VGND.n1561 VGND.n178 585
R320 VGND.n178 VGND.n97 585
R321 VGND.n1561 VGND.n190 585
R322 VGND.n190 VGND.n97 585
R323 VGND.n1561 VGND.n177 585
R324 VGND.n177 VGND.n97 585
R325 VGND.n1561 VGND.n193 585
R326 VGND.n193 VGND.n97 585
R327 VGND.n1561 VGND.n176 585
R328 VGND.n176 VGND.n97 585
R329 VGND.n1561 VGND.n196 585
R330 VGND.n196 VGND.n97 585
R331 VGND.n1561 VGND.n175 585
R332 VGND.n175 VGND.n97 585
R333 VGND.n1561 VGND.n199 585
R334 VGND.n199 VGND.n97 585
R335 VGND.n1561 VGND.n174 585
R336 VGND.n174 VGND.n97 585
R337 VGND.n1561 VGND.n202 585
R338 VGND.n202 VGND.n97 585
R339 VGND.n1561 VGND.n173 585
R340 VGND.n173 VGND.n97 585
R341 VGND.n1561 VGND.n205 585
R342 VGND.n205 VGND.n97 585
R343 VGND.n1561 VGND.n172 585
R344 VGND.n172 VGND.n97 585
R345 VGND.n1561 VGND.n208 585
R346 VGND.n208 VGND.n97 585
R347 VGND.n1561 VGND.n171 585
R348 VGND.n171 VGND.n97 585
R349 VGND.n1561 VGND.n211 585
R350 VGND.n211 VGND.n97 585
R351 VGND.n1561 VGND.n170 585
R352 VGND.n170 VGND.n97 585
R353 VGND.n1561 VGND.n214 585
R354 VGND.n214 VGND.n97 585
R355 VGND.n1561 VGND.n169 585
R356 VGND.n169 VGND.n97 585
R357 VGND.n1561 VGND.n217 585
R358 VGND.n217 VGND.n97 585
R359 VGND.n1561 VGND.n168 585
R360 VGND.n168 VGND.n97 585
R361 VGND.n1561 VGND.n220 585
R362 VGND.n220 VGND.n97 585
R363 VGND.n1561 VGND.n167 585
R364 VGND.n167 VGND.n97 585
R365 VGND.n1561 VGND.n223 585
R366 VGND.n223 VGND.n97 585
R367 VGND.n1561 VGND.n166 585
R368 VGND.n166 VGND.n97 585
R369 VGND.n1561 VGND.n226 585
R370 VGND.n226 VGND.n97 585
R371 VGND.n1561 VGND.n165 585
R372 VGND.n165 VGND.n97 585
R373 VGND.n1561 VGND.n229 585
R374 VGND.n229 VGND.n97 585
R375 VGND.n1561 VGND.n164 585
R376 VGND.n164 VGND.n97 585
R377 VGND.n1561 VGND.n232 585
R378 VGND.n232 VGND.n97 585
R379 VGND.n1561 VGND.n163 585
R380 VGND.n163 VGND.n97 585
R381 VGND.n1561 VGND.n235 585
R382 VGND.n235 VGND.n97 585
R383 VGND.n1561 VGND.n162 585
R384 VGND.n162 VGND.n97 585
R385 VGND.n1561 VGND.n238 585
R386 VGND.n238 VGND.n97 585
R387 VGND.n1561 VGND.n161 585
R388 VGND.n161 VGND.n97 585
R389 VGND.n1561 VGND.n241 585
R390 VGND.n241 VGND.n97 585
R391 VGND.n1561 VGND.n160 585
R392 VGND.n160 VGND.n97 585
R393 VGND.n1561 VGND.n244 585
R394 VGND.n244 VGND.n97 585
R395 VGND.n1561 VGND.n159 585
R396 VGND.n159 VGND.n97 585
R397 VGND.n1561 VGND.n247 585
R398 VGND.n247 VGND.n97 585
R399 VGND.n1561 VGND.n158 585
R400 VGND.n158 VGND.n97 585
R401 VGND.n1561 VGND.n250 585
R402 VGND.n250 VGND.n97 585
R403 VGND.n1561 VGND.n157 585
R404 VGND.n157 VGND.n97 585
R405 VGND.n1561 VGND.n253 585
R406 VGND.n253 VGND.n97 585
R407 VGND.n1561 VGND.n156 585
R408 VGND.n156 VGND.n97 585
R409 VGND.n1561 VGND.n256 585
R410 VGND.n256 VGND.n97 585
R411 VGND.n1561 VGND.n155 585
R412 VGND.n155 VGND.n97 585
R413 VGND.n1561 VGND.n259 585
R414 VGND.n259 VGND.n97 585
R415 VGND.n1561 VGND.n154 585
R416 VGND.n154 VGND.n97 585
R417 VGND.n1561 VGND.n262 585
R418 VGND.n262 VGND.n97 585
R419 VGND.n1561 VGND.n153 585
R420 VGND.n153 VGND.n97 585
R421 VGND.n1561 VGND.n265 585
R422 VGND.n265 VGND.n97 585
R423 VGND.n1561 VGND.n152 585
R424 VGND.n152 VGND.n97 585
R425 VGND.n1561 VGND.n268 585
R426 VGND.n268 VGND.n97 585
R427 VGND.n1561 VGND.n151 585
R428 VGND.n151 VGND.n97 585
R429 VGND.n1561 VGND.n271 585
R430 VGND.n271 VGND.n97 585
R431 VGND.n1561 VGND.n150 585
R432 VGND.n150 VGND.n97 585
R433 VGND.n1561 VGND.n274 585
R434 VGND.n274 VGND.n97 585
R435 VGND.n1561 VGND.n149 585
R436 VGND.n149 VGND.n97 585
R437 VGND.n1561 VGND.n277 585
R438 VGND.n277 VGND.n97 585
R439 VGND.n1561 VGND.n148 585
R440 VGND.n148 VGND.n97 585
R441 VGND.n1561 VGND.n280 585
R442 VGND.n280 VGND.n97 585
R443 VGND.n1561 VGND.n147 585
R444 VGND.n147 VGND.n97 585
R445 VGND.n1561 VGND.n283 585
R446 VGND.n283 VGND.n97 585
R447 VGND.n1561 VGND.n146 585
R448 VGND.n146 VGND.n97 585
R449 VGND.n1561 VGND.n286 585
R450 VGND.n286 VGND.n97 585
R451 VGND.n1561 VGND.n145 585
R452 VGND.n145 VGND.n97 585
R453 VGND.n1561 VGND.n289 585
R454 VGND.n289 VGND.n97 585
R455 VGND.n1561 VGND.n144 585
R456 VGND.n144 VGND.n97 585
R457 VGND.n1561 VGND.n292 585
R458 VGND.n292 VGND.n97 585
R459 VGND.n1561 VGND.n143 585
R460 VGND.n143 VGND.n97 585
R461 VGND.n1561 VGND.n295 585
R462 VGND.n295 VGND.n97 585
R463 VGND.n1561 VGND.n142 585
R464 VGND.n142 VGND.n97 585
R465 VGND.n1561 VGND.n298 585
R466 VGND.n298 VGND.n97 585
R467 VGND.n1561 VGND.n141 585
R468 VGND.n141 VGND.n97 585
R469 VGND.n1561 VGND.n301 585
R470 VGND.n301 VGND.n97 585
R471 VGND.n1561 VGND.n140 585
R472 VGND.n140 VGND.n97 585
R473 VGND.n1561 VGND.n304 585
R474 VGND.n304 VGND.n97 585
R475 VGND.n1561 VGND.n139 585
R476 VGND.n139 VGND.n97 585
R477 VGND.n1561 VGND.n307 585
R478 VGND.n307 VGND.n97 585
R479 VGND.n1561 VGND.n138 585
R480 VGND.n138 VGND.n97 585
R481 VGND.n1561 VGND.n310 585
R482 VGND.n310 VGND.n97 585
R483 VGND.n1561 VGND.n137 585
R484 VGND.n137 VGND.n97 585
R485 VGND.n1561 VGND.n313 585
R486 VGND.n313 VGND.n97 585
R487 VGND.n1561 VGND.n136 585
R488 VGND.n136 VGND.n97 585
R489 VGND.n1561 VGND.n316 585
R490 VGND.n316 VGND.n97 585
R491 VGND.n1561 VGND.n135 585
R492 VGND.n135 VGND.n97 585
R493 VGND.n1561 VGND.n319 585
R494 VGND.n319 VGND.n97 585
R495 VGND.n1561 VGND.n134 585
R496 VGND.n134 VGND.n97 585
R497 VGND.n1561 VGND.n322 585
R498 VGND.n322 VGND.n97 585
R499 VGND.n1561 VGND.n133 585
R500 VGND.n133 VGND.n97 585
R501 VGND.n1561 VGND.n325 585
R502 VGND.n325 VGND.n97 585
R503 VGND.n1561 VGND.n132 585
R504 VGND.n132 VGND.n97 585
R505 VGND.n1561 VGND.n328 585
R506 VGND.n328 VGND.n97 585
R507 VGND.n1561 VGND.n131 585
R508 VGND.n131 VGND.n97 585
R509 VGND.n1561 VGND.n331 585
R510 VGND.n331 VGND.n97 585
R511 VGND.n1561 VGND.n130 585
R512 VGND.n130 VGND.n97 585
R513 VGND.n1561 VGND.n334 585
R514 VGND.n334 VGND.n97 585
R515 VGND.n1561 VGND.n129 585
R516 VGND.n129 VGND.n97 585
R517 VGND.n1561 VGND.n337 585
R518 VGND.n337 VGND.n97 585
R519 VGND.n1561 VGND.n128 585
R520 VGND.n128 VGND.n97 585
R521 VGND.n1561 VGND.n340 585
R522 VGND.n340 VGND.n97 585
R523 VGND.n1561 VGND.n127 585
R524 VGND.n127 VGND.n97 585
R525 VGND.n1561 VGND.n343 585
R526 VGND.n343 VGND.n97 585
R527 VGND.n1561 VGND.n126 585
R528 VGND.n126 VGND.n97 585
R529 VGND.n1561 VGND.n346 585
R530 VGND.n346 VGND.n97 585
R531 VGND.n1561 VGND.n125 585
R532 VGND.n125 VGND.n97 585
R533 VGND.n1561 VGND.n349 585
R534 VGND.n349 VGND.n97 585
R535 VGND.n1561 VGND.n124 585
R536 VGND.n124 VGND.n97 585
R537 VGND.n1561 VGND.n352 585
R538 VGND.n352 VGND.n97 585
R539 VGND.n1561 VGND.n123 585
R540 VGND.n123 VGND.n97 585
R541 VGND.n1561 VGND.n355 585
R542 VGND.n355 VGND.n97 585
R543 VGND.n1561 VGND.n122 585
R544 VGND.n122 VGND.n97 585
R545 VGND.n1561 VGND.n358 585
R546 VGND.n358 VGND.n97 585
R547 VGND.n1561 VGND.n121 585
R548 VGND.n121 VGND.n97 585
R549 VGND.n1561 VGND.n361 585
R550 VGND.n361 VGND.n97 585
R551 VGND.n1561 VGND.n120 585
R552 VGND.n120 VGND.n97 585
R553 VGND.n1561 VGND.n364 585
R554 VGND.n364 VGND.n97 585
R555 VGND.n1561 VGND.n119 585
R556 VGND.n119 VGND.n97 585
R557 VGND.n1561 VGND.n367 585
R558 VGND.n367 VGND.n97 585
R559 VGND.n1561 VGND.n118 585
R560 VGND.n118 VGND.n97 585
R561 VGND.n1561 VGND.n370 585
R562 VGND.n370 VGND.n97 585
R563 VGND.n1561 VGND.n117 585
R564 VGND.n117 VGND.n97 585
R565 VGND.n1561 VGND.n373 585
R566 VGND.n373 VGND.n97 585
R567 VGND.n1561 VGND.n116 585
R568 VGND.n116 VGND.n97 585
R569 VGND.n1561 VGND.n376 585
R570 VGND.n376 VGND.n97 585
R571 VGND.n1561 VGND.n115 585
R572 VGND.n115 VGND.n97 585
R573 VGND.n1561 VGND.n379 585
R574 VGND.n379 VGND.n97 585
R575 VGND.n1561 VGND.n114 585
R576 VGND.n114 VGND.n97 585
R577 VGND.n1561 VGND.n382 585
R578 VGND.n382 VGND.n97 585
R579 VGND.n1561 VGND.n113 585
R580 VGND.n113 VGND.n97 585
R581 VGND.n1561 VGND.n385 585
R582 VGND.n385 VGND.n97 585
R583 VGND.n1561 VGND.n112 585
R584 VGND.n112 VGND.n97 585
R585 VGND.n1561 VGND.n388 585
R586 VGND.n388 VGND.n97 585
R587 VGND.n1561 VGND.n111 585
R588 VGND.n111 VGND.n97 585
R589 VGND.n1561 VGND.n391 585
R590 VGND.n391 VGND.n97 585
R591 VGND.n1561 VGND.n110 585
R592 VGND.n110 VGND.n97 585
R593 VGND.n1561 VGND.n394 585
R594 VGND.n394 VGND.n97 585
R595 VGND.n1561 VGND.n109 585
R596 VGND.n109 VGND.n97 585
R597 VGND.n1561 VGND.n397 585
R598 VGND.n397 VGND.n97 585
R599 VGND.n1561 VGND.n108 585
R600 VGND.n108 VGND.n97 585
R601 VGND.n1561 VGND.n400 585
R602 VGND.n400 VGND.n97 585
R603 VGND.n1561 VGND.n107 585
R604 VGND.n107 VGND.n97 585
R605 VGND.n1561 VGND.n403 585
R606 VGND.n403 VGND.n97 585
R607 VGND.n1561 VGND.n106 585
R608 VGND.n106 VGND.n97 585
R609 VGND.n1561 VGND.n406 585
R610 VGND.n406 VGND.n97 585
R611 VGND.n1561 VGND.n105 585
R612 VGND.n105 VGND.n97 585
R613 VGND.n1561 VGND.n1560 585
R614 VGND.n1560 VGND.n97 585
R615 VGND.n1561 VGND.n104 585
R616 VGND.n104 VGND.n97 585
R617 VGND.n1562 VGND.n103 585
R618 VGND.n1562 VGND.n1561 585
R619 VGND.n1562 VGND.n97 585
R620 VGND.n859 VGND.n626 281.14
R621 VGND.n939 VGND.n938 281.14
R622 VGND.n857 VGND.n626 281.14
R623 VGND.n938 VGND.n862 281.14
R624 VGND.n855 VGND.n626 281.14
R625 VGND.n938 VGND.n863 281.14
R626 VGND.n853 VGND.n626 281.14
R627 VGND.n938 VGND.n864 281.14
R628 VGND.n851 VGND.n626 281.14
R629 VGND.n938 VGND.n865 281.14
R630 VGND.n849 VGND.n626 281.14
R631 VGND.n938 VGND.n866 281.14
R632 VGND.n847 VGND.n626 281.14
R633 VGND.n938 VGND.n867 281.14
R634 VGND.n845 VGND.n626 281.14
R635 VGND.n938 VGND.n868 281.14
R636 VGND.n843 VGND.n626 281.14
R637 VGND.n938 VGND.n869 281.14
R638 VGND.n841 VGND.n626 281.14
R639 VGND.n938 VGND.n870 281.14
R640 VGND.n839 VGND.n626 281.14
R641 VGND.n938 VGND.n871 281.14
R642 VGND.n837 VGND.n626 281.14
R643 VGND.n938 VGND.n872 281.14
R644 VGND.n835 VGND.n626 281.14
R645 VGND.n938 VGND.n873 281.14
R646 VGND.n833 VGND.n626 281.14
R647 VGND.n938 VGND.n874 281.14
R648 VGND.n831 VGND.n626 281.14
R649 VGND.n938 VGND.n875 281.14
R650 VGND.n829 VGND.n626 281.14
R651 VGND.n938 VGND.n876 281.14
R652 VGND.n827 VGND.n626 281.14
R653 VGND.n938 VGND.n877 281.14
R654 VGND.n825 VGND.n626 281.14
R655 VGND.n938 VGND.n878 281.14
R656 VGND.n823 VGND.n626 281.14
R657 VGND.n938 VGND.n879 281.14
R658 VGND.n821 VGND.n626 281.14
R659 VGND.n938 VGND.n880 281.14
R660 VGND.n819 VGND.n626 281.14
R661 VGND.n938 VGND.n881 281.14
R662 VGND.n817 VGND.n626 281.14
R663 VGND.n938 VGND.n882 281.14
R664 VGND.n815 VGND.n626 281.14
R665 VGND.n938 VGND.n883 281.14
R666 VGND.n813 VGND.n626 281.14
R667 VGND.n938 VGND.n884 281.14
R668 VGND.n811 VGND.n626 281.14
R669 VGND.n938 VGND.n885 281.14
R670 VGND.n809 VGND.n626 281.14
R671 VGND.n938 VGND.n886 281.14
R672 VGND.n807 VGND.n626 281.14
R673 VGND.n938 VGND.n887 281.14
R674 VGND.n805 VGND.n626 281.14
R675 VGND.n938 VGND.n888 281.14
R676 VGND.n803 VGND.n626 281.14
R677 VGND.n938 VGND.n889 281.14
R678 VGND.n801 VGND.n626 281.14
R679 VGND.n938 VGND.n890 281.14
R680 VGND.n799 VGND.n626 281.14
R681 VGND.n938 VGND.n891 281.14
R682 VGND.n797 VGND.n626 281.14
R683 VGND.n938 VGND.n892 281.14
R684 VGND.n795 VGND.n626 281.14
R685 VGND.n938 VGND.n893 281.14
R686 VGND.n793 VGND.n626 281.14
R687 VGND.n938 VGND.n894 281.14
R688 VGND.n791 VGND.n626 281.14
R689 VGND.n938 VGND.n895 281.14
R690 VGND.n789 VGND.n626 281.14
R691 VGND.n938 VGND.n896 281.14
R692 VGND.n787 VGND.n626 281.14
R693 VGND.n938 VGND.n897 281.14
R694 VGND.n785 VGND.n626 281.14
R695 VGND.n938 VGND.n898 281.14
R696 VGND.n783 VGND.n626 281.14
R697 VGND.n938 VGND.n899 281.14
R698 VGND.n781 VGND.n626 281.14
R699 VGND.n938 VGND.n900 281.14
R700 VGND.n779 VGND.n626 281.14
R701 VGND.n938 VGND.n901 281.14
R702 VGND.n777 VGND.n626 281.14
R703 VGND.n938 VGND.n902 281.14
R704 VGND.n775 VGND.n626 281.14
R705 VGND.n938 VGND.n903 281.14
R706 VGND.n773 VGND.n626 281.14
R707 VGND.n938 VGND.n904 281.14
R708 VGND.n771 VGND.n626 281.14
R709 VGND.n938 VGND.n905 281.14
R710 VGND.n769 VGND.n626 281.14
R711 VGND.n938 VGND.n906 281.14
R712 VGND.n767 VGND.n626 281.14
R713 VGND.n938 VGND.n907 281.14
R714 VGND.n765 VGND.n626 281.14
R715 VGND.n938 VGND.n908 281.14
R716 VGND.n763 VGND.n626 281.14
R717 VGND.n938 VGND.n909 281.14
R718 VGND.n761 VGND.n626 281.14
R719 VGND.n938 VGND.n910 281.14
R720 VGND.n759 VGND.n626 281.14
R721 VGND.n938 VGND.n911 281.14
R722 VGND.n757 VGND.n626 281.14
R723 VGND.n938 VGND.n912 281.14
R724 VGND.n755 VGND.n626 281.14
R725 VGND.n938 VGND.n913 281.14
R726 VGND.n753 VGND.n626 281.14
R727 VGND.n938 VGND.n914 281.14
R728 VGND.n751 VGND.n626 281.14
R729 VGND.n938 VGND.n915 281.14
R730 VGND.n749 VGND.n626 281.14
R731 VGND.n938 VGND.n916 281.14
R732 VGND.n747 VGND.n626 281.14
R733 VGND.n938 VGND.n917 281.14
R734 VGND.n745 VGND.n626 281.14
R735 VGND.n938 VGND.n918 281.14
R736 VGND.n743 VGND.n626 281.14
R737 VGND.n938 VGND.n919 281.14
R738 VGND.n741 VGND.n626 281.14
R739 VGND.n938 VGND.n920 281.14
R740 VGND.n739 VGND.n626 281.14
R741 VGND.n938 VGND.n921 281.14
R742 VGND.n737 VGND.n626 281.14
R743 VGND.n938 VGND.n922 281.14
R744 VGND.n735 VGND.n626 281.14
R745 VGND.n938 VGND.n923 281.14
R746 VGND.n733 VGND.n626 281.14
R747 VGND.n938 VGND.n924 281.14
R748 VGND.n731 VGND.n626 281.14
R749 VGND.n938 VGND.n925 281.14
R750 VGND.n729 VGND.n626 281.14
R751 VGND.n938 VGND.n926 281.14
R752 VGND.n727 VGND.n626 281.14
R753 VGND.n938 VGND.n927 281.14
R754 VGND.n725 VGND.n626 281.14
R755 VGND.n938 VGND.n928 281.14
R756 VGND.n723 VGND.n626 281.14
R757 VGND.n938 VGND.n929 281.14
R758 VGND.n721 VGND.n626 281.14
R759 VGND.n938 VGND.n930 281.14
R760 VGND.n719 VGND.n626 281.14
R761 VGND.n938 VGND.n931 281.14
R762 VGND.n717 VGND.n626 281.14
R763 VGND.n938 VGND.n932 281.14
R764 VGND.n715 VGND.n626 281.14
R765 VGND.n938 VGND.n933 281.14
R766 VGND.n713 VGND.n626 281.14
R767 VGND.n938 VGND.n934 281.14
R768 VGND.n711 VGND.n626 281.14
R769 VGND.n938 VGND.n935 281.14
R770 VGND.n709 VGND.n626 281.14
R771 VGND.n938 VGND.n936 281.14
R772 VGND.n938 VGND.n631 281.14
R773 VGND.n183 VGND.n96 281.14
R774 VGND.n182 VGND.n103 281.14
R775 VGND.n186 VGND.n96 281.14
R776 VGND.n185 VGND.n103 281.14
R777 VGND.n189 VGND.n96 281.14
R778 VGND.n188 VGND.n103 281.14
R779 VGND.n192 VGND.n96 281.14
R780 VGND.n191 VGND.n103 281.14
R781 VGND.n195 VGND.n96 281.14
R782 VGND.n194 VGND.n103 281.14
R783 VGND.n198 VGND.n96 281.14
R784 VGND.n197 VGND.n103 281.14
R785 VGND.n201 VGND.n96 281.14
R786 VGND.n200 VGND.n103 281.14
R787 VGND.n204 VGND.n96 281.14
R788 VGND.n203 VGND.n103 281.14
R789 VGND.n207 VGND.n96 281.14
R790 VGND.n206 VGND.n103 281.14
R791 VGND.n210 VGND.n96 281.14
R792 VGND.n209 VGND.n103 281.14
R793 VGND.n213 VGND.n96 281.14
R794 VGND.n212 VGND.n103 281.14
R795 VGND.n216 VGND.n96 281.14
R796 VGND.n215 VGND.n103 281.14
R797 VGND.n219 VGND.n96 281.14
R798 VGND.n218 VGND.n103 281.14
R799 VGND.n222 VGND.n96 281.14
R800 VGND.n221 VGND.n103 281.14
R801 VGND.n225 VGND.n96 281.14
R802 VGND.n224 VGND.n103 281.14
R803 VGND.n228 VGND.n96 281.14
R804 VGND.n227 VGND.n103 281.14
R805 VGND.n231 VGND.n96 281.14
R806 VGND.n230 VGND.n103 281.14
R807 VGND.n234 VGND.n96 281.14
R808 VGND.n233 VGND.n103 281.14
R809 VGND.n237 VGND.n96 281.14
R810 VGND.n236 VGND.n103 281.14
R811 VGND.n240 VGND.n96 281.14
R812 VGND.n239 VGND.n103 281.14
R813 VGND.n243 VGND.n96 281.14
R814 VGND.n242 VGND.n103 281.14
R815 VGND.n246 VGND.n96 281.14
R816 VGND.n245 VGND.n103 281.14
R817 VGND.n249 VGND.n96 281.14
R818 VGND.n248 VGND.n103 281.14
R819 VGND.n252 VGND.n96 281.14
R820 VGND.n251 VGND.n103 281.14
R821 VGND.n255 VGND.n96 281.14
R822 VGND.n254 VGND.n103 281.14
R823 VGND.n258 VGND.n96 281.14
R824 VGND.n257 VGND.n103 281.14
R825 VGND.n261 VGND.n96 281.14
R826 VGND.n260 VGND.n103 281.14
R827 VGND.n264 VGND.n96 281.14
R828 VGND.n263 VGND.n103 281.14
R829 VGND.n267 VGND.n96 281.14
R830 VGND.n266 VGND.n103 281.14
R831 VGND.n270 VGND.n96 281.14
R832 VGND.n269 VGND.n103 281.14
R833 VGND.n273 VGND.n96 281.14
R834 VGND.n272 VGND.n103 281.14
R835 VGND.n276 VGND.n96 281.14
R836 VGND.n275 VGND.n103 281.14
R837 VGND.n279 VGND.n96 281.14
R838 VGND.n278 VGND.n103 281.14
R839 VGND.n282 VGND.n96 281.14
R840 VGND.n281 VGND.n103 281.14
R841 VGND.n285 VGND.n96 281.14
R842 VGND.n284 VGND.n103 281.14
R843 VGND.n288 VGND.n96 281.14
R844 VGND.n287 VGND.n103 281.14
R845 VGND.n291 VGND.n96 281.14
R846 VGND.n290 VGND.n103 281.14
R847 VGND.n294 VGND.n96 281.14
R848 VGND.n293 VGND.n103 281.14
R849 VGND.n297 VGND.n96 281.14
R850 VGND.n296 VGND.n103 281.14
R851 VGND.n300 VGND.n96 281.14
R852 VGND.n299 VGND.n103 281.14
R853 VGND.n303 VGND.n96 281.14
R854 VGND.n302 VGND.n103 281.14
R855 VGND.n306 VGND.n96 281.14
R856 VGND.n305 VGND.n103 281.14
R857 VGND.n309 VGND.n96 281.14
R858 VGND.n308 VGND.n103 281.14
R859 VGND.n312 VGND.n96 281.14
R860 VGND.n311 VGND.n103 281.14
R861 VGND.n315 VGND.n96 281.14
R862 VGND.n314 VGND.n103 281.14
R863 VGND.n318 VGND.n96 281.14
R864 VGND.n317 VGND.n103 281.14
R865 VGND.n321 VGND.n96 281.14
R866 VGND.n320 VGND.n103 281.14
R867 VGND.n324 VGND.n96 281.14
R868 VGND.n323 VGND.n103 281.14
R869 VGND.n327 VGND.n96 281.14
R870 VGND.n326 VGND.n103 281.14
R871 VGND.n330 VGND.n96 281.14
R872 VGND.n329 VGND.n103 281.14
R873 VGND.n333 VGND.n96 281.14
R874 VGND.n332 VGND.n103 281.14
R875 VGND.n336 VGND.n96 281.14
R876 VGND.n335 VGND.n103 281.14
R877 VGND.n339 VGND.n96 281.14
R878 VGND.n338 VGND.n103 281.14
R879 VGND.n342 VGND.n96 281.14
R880 VGND.n341 VGND.n103 281.14
R881 VGND.n345 VGND.n96 281.14
R882 VGND.n344 VGND.n103 281.14
R883 VGND.n348 VGND.n96 281.14
R884 VGND.n347 VGND.n103 281.14
R885 VGND.n351 VGND.n96 281.14
R886 VGND.n350 VGND.n103 281.14
R887 VGND.n354 VGND.n96 281.14
R888 VGND.n353 VGND.n103 281.14
R889 VGND.n357 VGND.n96 281.14
R890 VGND.n356 VGND.n103 281.14
R891 VGND.n360 VGND.n96 281.14
R892 VGND.n359 VGND.n103 281.14
R893 VGND.n363 VGND.n96 281.14
R894 VGND.n362 VGND.n103 281.14
R895 VGND.n366 VGND.n96 281.14
R896 VGND.n365 VGND.n103 281.14
R897 VGND.n369 VGND.n96 281.14
R898 VGND.n368 VGND.n103 281.14
R899 VGND.n372 VGND.n96 281.14
R900 VGND.n371 VGND.n103 281.14
R901 VGND.n375 VGND.n96 281.14
R902 VGND.n374 VGND.n103 281.14
R903 VGND.n378 VGND.n96 281.14
R904 VGND.n377 VGND.n103 281.14
R905 VGND.n381 VGND.n96 281.14
R906 VGND.n380 VGND.n103 281.14
R907 VGND.n384 VGND.n96 281.14
R908 VGND.n383 VGND.n103 281.14
R909 VGND.n387 VGND.n96 281.14
R910 VGND.n386 VGND.n103 281.14
R911 VGND.n390 VGND.n96 281.14
R912 VGND.n389 VGND.n103 281.14
R913 VGND.n393 VGND.n96 281.14
R914 VGND.n392 VGND.n103 281.14
R915 VGND.n396 VGND.n96 281.14
R916 VGND.n395 VGND.n103 281.14
R917 VGND.n399 VGND.n96 281.14
R918 VGND.n398 VGND.n103 281.14
R919 VGND.n402 VGND.n96 281.14
R920 VGND.n401 VGND.n103 281.14
R921 VGND.n405 VGND.n96 281.14
R922 VGND.n404 VGND.n103 281.14
R923 VGND.n408 VGND.n96 281.14
R924 VGND.n407 VGND.n103 281.14
R925 VGND.n102 VGND.n96 281.14
R926 VGND.n941 VGND.n629 166.845
R927 VGND.n1567 VGND.n1566 166.845
R928 VGND.n1566 VGND.n1565 166.843
R929 VGND.n1103 VGND.n629 166.843
R930 VGND.n1098 VGND.n1097 146.25
R931 VGND.n1096 VGND.n633 146.25
R932 VGND.n1095 VGND.n860 146.25
R933 VGND.n1094 VGND.n634 146.25
R934 VGND.n1093 VGND.n858 146.25
R935 VGND.n1092 VGND.n635 146.25
R936 VGND.n1091 VGND.n856 146.25
R937 VGND.n1090 VGND.n636 146.25
R938 VGND.n1089 VGND.n854 146.25
R939 VGND.n1088 VGND.n637 146.25
R940 VGND.n1087 VGND.n852 146.25
R941 VGND.n1086 VGND.n638 146.25
R942 VGND.n1085 VGND.n850 146.25
R943 VGND.n1084 VGND.n639 146.25
R944 VGND.n1083 VGND.n848 146.25
R945 VGND.n1082 VGND.n640 146.25
R946 VGND.n1081 VGND.n846 146.25
R947 VGND.n1080 VGND.n641 146.25
R948 VGND.n1079 VGND.n844 146.25
R949 VGND.n1078 VGND.n642 146.25
R950 VGND.n1077 VGND.n842 146.25
R951 VGND.n1076 VGND.n643 146.25
R952 VGND.n1075 VGND.n840 146.25
R953 VGND.n1074 VGND.n644 146.25
R954 VGND.n1073 VGND.n838 146.25
R955 VGND.n1072 VGND.n645 146.25
R956 VGND.n1071 VGND.n836 146.25
R957 VGND.n1070 VGND.n646 146.25
R958 VGND.n1069 VGND.n834 146.25
R959 VGND.n1068 VGND.n647 146.25
R960 VGND.n1067 VGND.n832 146.25
R961 VGND.n1066 VGND.n648 146.25
R962 VGND.n1065 VGND.n830 146.25
R963 VGND.n1064 VGND.n649 146.25
R964 VGND.n1063 VGND.n828 146.25
R965 VGND.n1062 VGND.n650 146.25
R966 VGND.n1061 VGND.n826 146.25
R967 VGND.n1060 VGND.n651 146.25
R968 VGND.n1059 VGND.n824 146.25
R969 VGND.n1058 VGND.n652 146.25
R970 VGND.n1057 VGND.n822 146.25
R971 VGND.n1056 VGND.n653 146.25
R972 VGND.n1055 VGND.n820 146.25
R973 VGND.n1054 VGND.n654 146.25
R974 VGND.n1053 VGND.n818 146.25
R975 VGND.n1052 VGND.n655 146.25
R976 VGND.n1051 VGND.n816 146.25
R977 VGND.n1050 VGND.n656 146.25
R978 VGND.n1049 VGND.n814 146.25
R979 VGND.n1048 VGND.n657 146.25
R980 VGND.n1047 VGND.n812 146.25
R981 VGND.n1046 VGND.n658 146.25
R982 VGND.n1045 VGND.n810 146.25
R983 VGND.n1044 VGND.n659 146.25
R984 VGND.n1043 VGND.n808 146.25
R985 VGND.n1042 VGND.n660 146.25
R986 VGND.n1041 VGND.n806 146.25
R987 VGND.n1040 VGND.n661 146.25
R988 VGND.n1039 VGND.n804 146.25
R989 VGND.n1038 VGND.n662 146.25
R990 VGND.n1037 VGND.n802 146.25
R991 VGND.n1036 VGND.n663 146.25
R992 VGND.n1035 VGND.n800 146.25
R993 VGND.n1034 VGND.n664 146.25
R994 VGND.n1033 VGND.n798 146.25
R995 VGND.n1032 VGND.n665 146.25
R996 VGND.n1031 VGND.n796 146.25
R997 VGND.n1030 VGND.n666 146.25
R998 VGND.n1029 VGND.n794 146.25
R999 VGND.n1028 VGND.n667 146.25
R1000 VGND.n1027 VGND.n792 146.25
R1001 VGND.n1026 VGND.n668 146.25
R1002 VGND.n1025 VGND.n790 146.25
R1003 VGND.n1024 VGND.n669 146.25
R1004 VGND.n1023 VGND.n788 146.25
R1005 VGND.n1022 VGND.n670 146.25
R1006 VGND.n1021 VGND.n786 146.25
R1007 VGND.n1018 VGND.n671 146.25
R1008 VGND.n1017 VGND.n784 146.25
R1009 VGND.n1016 VGND.n672 146.25
R1010 VGND.n1015 VGND.n782 146.25
R1011 VGND.n1014 VGND.n673 146.25
R1012 VGND.n1013 VGND.n780 146.25
R1013 VGND.n1012 VGND.n674 146.25
R1014 VGND.n1011 VGND.n778 146.25
R1015 VGND.n1010 VGND.n675 146.25
R1016 VGND.n1009 VGND.n776 146.25
R1017 VGND.n1008 VGND.n676 146.25
R1018 VGND.n1007 VGND.n774 146.25
R1019 VGND.n1006 VGND.n677 146.25
R1020 VGND.n1005 VGND.n772 146.25
R1021 VGND.n1004 VGND.n678 146.25
R1022 VGND.n1003 VGND.n770 146.25
R1023 VGND.n1002 VGND.n679 146.25
R1024 VGND.n1001 VGND.n768 146.25
R1025 VGND.n1000 VGND.n680 146.25
R1026 VGND.n999 VGND.n766 146.25
R1027 VGND.n998 VGND.n681 146.25
R1028 VGND.n997 VGND.n764 146.25
R1029 VGND.n996 VGND.n682 146.25
R1030 VGND.n995 VGND.n762 146.25
R1031 VGND.n994 VGND.n683 146.25
R1032 VGND.n993 VGND.n760 146.25
R1033 VGND.n992 VGND.n684 146.25
R1034 VGND.n991 VGND.n758 146.25
R1035 VGND.n990 VGND.n685 146.25
R1036 VGND.n989 VGND.n756 146.25
R1037 VGND.n988 VGND.n686 146.25
R1038 VGND.n987 VGND.n754 146.25
R1039 VGND.n986 VGND.n687 146.25
R1040 VGND.n985 VGND.n752 146.25
R1041 VGND.n984 VGND.n688 146.25
R1042 VGND.n983 VGND.n750 146.25
R1043 VGND.n982 VGND.n689 146.25
R1044 VGND.n981 VGND.n748 146.25
R1045 VGND.n980 VGND.n690 146.25
R1046 VGND.n979 VGND.n746 146.25
R1047 VGND.n978 VGND.n691 146.25
R1048 VGND.n977 VGND.n744 146.25
R1049 VGND.n976 VGND.n692 146.25
R1050 VGND.n975 VGND.n742 146.25
R1051 VGND.n974 VGND.n693 146.25
R1052 VGND.n973 VGND.n740 146.25
R1053 VGND.n972 VGND.n694 146.25
R1054 VGND.n971 VGND.n738 146.25
R1055 VGND.n970 VGND.n695 146.25
R1056 VGND.n969 VGND.n736 146.25
R1057 VGND.n968 VGND.n696 146.25
R1058 VGND.n967 VGND.n734 146.25
R1059 VGND.n966 VGND.n697 146.25
R1060 VGND.n965 VGND.n732 146.25
R1061 VGND.n964 VGND.n698 146.25
R1062 VGND.n963 VGND.n730 146.25
R1063 VGND.n962 VGND.n699 146.25
R1064 VGND.n961 VGND.n728 146.25
R1065 VGND.n960 VGND.n700 146.25
R1066 VGND.n959 VGND.n726 146.25
R1067 VGND.n958 VGND.n701 146.25
R1068 VGND.n957 VGND.n724 146.25
R1069 VGND.n956 VGND.n702 146.25
R1070 VGND.n955 VGND.n722 146.25
R1071 VGND.n954 VGND.n703 146.25
R1072 VGND.n953 VGND.n720 146.25
R1073 VGND.n952 VGND.n704 146.25
R1074 VGND.n951 VGND.n718 146.25
R1075 VGND.n950 VGND.n705 146.25
R1076 VGND.n949 VGND.n716 146.25
R1077 VGND.n948 VGND.n706 146.25
R1078 VGND.n947 VGND.n714 146.25
R1079 VGND.n946 VGND.n707 146.25
R1080 VGND.n945 VGND.n712 146.25
R1081 VGND.n944 VGND.n708 146.25
R1082 VGND.n943 VGND.n710 146.25
R1083 VGND.n1100 VGND.n628 146.25
R1084 VGND.n940 VGND.n630 146.25
R1085 VGND.n625 VGND.n624 146.25
R1086 VGND.n937 VGND.n625 146.25
R1087 VGND.n1110 VGND.n1109 146.25
R1088 VGND.n1109 VGND.n1108 146.25
R1089 VGND.n1111 VGND.n623 146.25
R1090 VGND.n623 VGND.n622 146.25
R1091 VGND.n1113 VGND.n1112 146.25
R1092 VGND.n1114 VGND.n1113 146.25
R1093 VGND.n617 VGND.n616 146.25
R1094 VGND.n618 VGND.n617 146.25
R1095 VGND.n1122 VGND.n1121 146.25
R1096 VGND.n1121 VGND.n1120 146.25
R1097 VGND.n1123 VGND.n615 146.25
R1098 VGND.n615 VGND.n614 146.25
R1099 VGND.n1125 VGND.n1124 146.25
R1100 VGND.n1126 VGND.n1125 146.25
R1101 VGND.n608 VGND.n607 146.25
R1102 VGND.n609 VGND.n608 146.25
R1103 VGND.n1134 VGND.n1133 146.25
R1104 VGND.n1133 VGND.n1132 146.25
R1105 VGND.n1135 VGND.n606 146.25
R1106 VGND.n610 VGND.n606 146.25
R1107 VGND.n1137 VGND.n1136 146.25
R1108 VGND.n1138 VGND.n1137 146.25
R1109 VGND.n601 VGND.n600 146.25
R1110 VGND.n602 VGND.n601 146.25
R1111 VGND.n1146 VGND.n1145 146.25
R1112 VGND.n1145 VGND.n1144 146.25
R1113 VGND.n1147 VGND.n599 146.25
R1114 VGND.n599 VGND.n598 146.25
R1115 VGND.n1149 VGND.n1148 146.25
R1116 VGND.n1150 VGND.n1149 146.25
R1117 VGND.n593 VGND.n592 146.25
R1118 VGND.n594 VGND.n593 146.25
R1119 VGND.n1158 VGND.n1157 146.25
R1120 VGND.n1157 VGND.n1156 146.25
R1121 VGND.n1159 VGND.n591 146.25
R1122 VGND.n591 VGND.n589 146.25
R1123 VGND.n1161 VGND.n1160 146.25
R1124 VGND.n1162 VGND.n1161 146.25
R1125 VGND.n585 VGND.n584 146.25
R1126 VGND.n590 VGND.n585 146.25
R1127 VGND.n1170 VGND.n1169 146.25
R1128 VGND.n1169 VGND.n1168 146.25
R1129 VGND.n1171 VGND.n583 146.25
R1130 VGND.n583 VGND.n582 146.25
R1131 VGND.n1173 VGND.n1172 146.25
R1132 VGND.n1174 VGND.n1173 146.25
R1133 VGND.n577 VGND.n576 146.25
R1134 VGND.n578 VGND.n577 146.25
R1135 VGND.n1182 VGND.n1181 146.25
R1136 VGND.n1181 VGND.n1180 146.25
R1137 VGND.n1183 VGND.n575 146.25
R1138 VGND.n575 VGND.n574 146.25
R1139 VGND.n1185 VGND.n1184 146.25
R1140 VGND.n1186 VGND.n1185 146.25
R1141 VGND.n568 VGND.n567 146.25
R1142 VGND.n569 VGND.n568 146.25
R1143 VGND.n1194 VGND.n1193 146.25
R1144 VGND.n1193 VGND.n1192 146.25
R1145 VGND.n1195 VGND.n566 146.25
R1146 VGND.n570 VGND.n566 146.25
R1147 VGND.n1197 VGND.n1196 146.25
R1148 VGND.n1198 VGND.n1197 146.25
R1149 VGND.n561 VGND.n560 146.25
R1150 VGND.n562 VGND.n561 146.25
R1151 VGND.n1206 VGND.n1205 146.25
R1152 VGND.n1205 VGND.n1204 146.25
R1153 VGND.n1207 VGND.n559 146.25
R1154 VGND.n559 VGND.n558 146.25
R1155 VGND.n1209 VGND.n1208 146.25
R1156 VGND.n1210 VGND.n1209 146.25
R1157 VGND.n553 VGND.n552 146.25
R1158 VGND.n554 VGND.n553 146.25
R1159 VGND.n1218 VGND.n1217 146.25
R1160 VGND.n1217 VGND.n1216 146.25
R1161 VGND.n1219 VGND.n551 146.25
R1162 VGND.n551 VGND.n549 146.25
R1163 VGND.n1221 VGND.n1220 146.25
R1164 VGND.n1222 VGND.n1221 146.25
R1165 VGND.n545 VGND.n544 146.25
R1166 VGND.n550 VGND.n545 146.25
R1167 VGND.n1230 VGND.n1229 146.25
R1168 VGND.n1229 VGND.n1228 146.25
R1169 VGND.n1231 VGND.n543 146.25
R1170 VGND.n543 VGND.n542 146.25
R1171 VGND.n1233 VGND.n1232 146.25
R1172 VGND.n1234 VGND.n1233 146.25
R1173 VGND.n537 VGND.n536 146.25
R1174 VGND.n538 VGND.n537 146.25
R1175 VGND.n1242 VGND.n1241 146.25
R1176 VGND.n1241 VGND.n1240 146.25
R1177 VGND.n1243 VGND.n535 146.25
R1178 VGND.n535 VGND.n534 146.25
R1179 VGND.n1245 VGND.n1244 146.25
R1180 VGND.n1246 VGND.n1245 146.25
R1181 VGND.n528 VGND.n527 146.25
R1182 VGND.n529 VGND.n528 146.25
R1183 VGND.n1254 VGND.n1253 146.25
R1184 VGND.n1253 VGND.n1252 146.25
R1185 VGND.n1255 VGND.n526 146.25
R1186 VGND.n530 VGND.n526 146.25
R1187 VGND.n1257 VGND.n1256 146.25
R1188 VGND.n1258 VGND.n1257 146.25
R1189 VGND.n521 VGND.n520 146.25
R1190 VGND.n522 VGND.n521 146.25
R1191 VGND.n1266 VGND.n1265 146.25
R1192 VGND.n1265 VGND.n1264 146.25
R1193 VGND.n1267 VGND.n519 146.25
R1194 VGND.n519 VGND.n518 146.25
R1195 VGND.n1269 VGND.n1268 146.25
R1196 VGND.n1270 VGND.n1269 146.25
R1197 VGND.n513 VGND.n512 146.25
R1198 VGND.n514 VGND.n513 146.25
R1199 VGND.n1278 VGND.n1277 146.25
R1200 VGND.n1277 VGND.n1276 146.25
R1201 VGND.n1279 VGND.n511 146.25
R1202 VGND.n511 VGND.n509 146.25
R1203 VGND.n1281 VGND.n1280 146.25
R1204 VGND.n1282 VGND.n1281 146.25
R1205 VGND.n505 VGND.n504 146.25
R1206 VGND.n510 VGND.n505 146.25
R1207 VGND.n1290 VGND.n1289 146.25
R1208 VGND.n1289 VGND.n1288 146.25
R1209 VGND.n1291 VGND.n503 146.25
R1210 VGND.n503 VGND.n502 146.25
R1211 VGND.n1293 VGND.n1292 146.25
R1212 VGND.n1294 VGND.n1293 146.25
R1213 VGND.n497 VGND.n496 146.25
R1214 VGND.n498 VGND.n497 146.25
R1215 VGND.n1302 VGND.n1301 146.25
R1216 VGND.n1301 VGND.n1300 146.25
R1217 VGND.n1303 VGND.n494 146.25
R1218 VGND.n494 VGND.n492 146.25
R1219 VGND.n1308 VGND.n1307 146.25
R1220 VGND.n1309 VGND.n1308 146.25
R1221 VGND.n1306 VGND.n495 146.25
R1222 VGND.n495 VGND.n493 146.25
R1223 VGND.n1305 VGND.n1304 146.25
R1224 VGND.n1304 VGND.n488 146.25
R1225 VGND.n487 VGND.n486 146.25
R1226 VGND.n1316 VGND.n487 146.25
R1227 VGND.n1476 VGND.n1317 146.25
R1228 VGND.n1317 VGND.t15 146.25
R1229 VGND.n1475 VGND.n1474 146.25
R1230 VGND.n1474 VGND.n5 146.25
R1231 VGND.n1473 VGND.n1318 146.25
R1232 VGND.n1473 VGND.n6 146.25
R1233 VGND.n1472 VGND.n1471 146.25
R1234 VGND.n1472 VGND.n7 146.25
R1235 VGND.n1470 VGND.n1320 146.25
R1236 VGND.n1320 VGND.n1319 146.25
R1237 VGND.n1469 VGND.n1468 146.25
R1238 VGND.n1468 VGND.n10 146.25
R1239 VGND.n1467 VGND.n1321 146.25
R1240 VGND.n1467 VGND.n11 146.25
R1241 VGND.n1466 VGND.n1465 146.25
R1242 VGND.n1466 VGND.n12 146.25
R1243 VGND.n1464 VGND.n1323 146.25
R1244 VGND.n1323 VGND.n1322 146.25
R1245 VGND.n1463 VGND.n1462 146.25
R1246 VGND.n1462 VGND.n15 146.25
R1247 VGND.n1461 VGND.n1324 146.25
R1248 VGND.n1461 VGND.n16 146.25
R1249 VGND.n1460 VGND.n1459 146.25
R1250 VGND.n1460 VGND.n17 146.25
R1251 VGND.n1458 VGND.n1326 146.25
R1252 VGND.n1326 VGND.n1325 146.25
R1253 VGND.n1457 VGND.n1456 146.25
R1254 VGND.n1456 VGND.n20 146.25
R1255 VGND.n1455 VGND.n1327 146.25
R1256 VGND.n1455 VGND.n21 146.25
R1257 VGND.n1454 VGND.n1453 146.25
R1258 VGND.n1454 VGND.n22 146.25
R1259 VGND.n1452 VGND.n1329 146.25
R1260 VGND.n1329 VGND.n1328 146.25
R1261 VGND.n1451 VGND.n1450 146.25
R1262 VGND.n1450 VGND.n25 146.25
R1263 VGND.n1449 VGND.n1330 146.25
R1264 VGND.n1449 VGND.n26 146.25
R1265 VGND.n1448 VGND.n1447 146.25
R1266 VGND.n1448 VGND.n27 146.25
R1267 VGND.n1446 VGND.n1332 146.25
R1268 VGND.n1332 VGND.n1331 146.25
R1269 VGND.n1445 VGND.n1444 146.25
R1270 VGND.n1444 VGND.n30 146.25
R1271 VGND.n1443 VGND.n1333 146.25
R1272 VGND.n1443 VGND.n31 146.25
R1273 VGND.n1442 VGND.n1441 146.25
R1274 VGND.n1442 VGND.n32 146.25
R1275 VGND.n1440 VGND.n1335 146.25
R1276 VGND.n1335 VGND.n1334 146.25
R1277 VGND.n1439 VGND.n1438 146.25
R1278 VGND.n1438 VGND.n35 146.25
R1279 VGND.n1437 VGND.n1336 146.25
R1280 VGND.n1437 VGND.n36 146.25
R1281 VGND.n1436 VGND.n1435 146.25
R1282 VGND.n1436 VGND.n37 146.25
R1283 VGND.n1434 VGND.n1338 146.25
R1284 VGND.n1338 VGND.n1337 146.25
R1285 VGND.n1433 VGND.n1432 146.25
R1286 VGND.n1432 VGND.n40 146.25
R1287 VGND.n1431 VGND.n1339 146.25
R1288 VGND.n1431 VGND.n41 146.25
R1289 VGND.n1430 VGND.n1429 146.25
R1290 VGND.n1430 VGND.n42 146.25
R1291 VGND.n1428 VGND.n1341 146.25
R1292 VGND.n1341 VGND.n1340 146.25
R1293 VGND.n1427 VGND.n1426 146.25
R1294 VGND.n1426 VGND.n45 146.25
R1295 VGND.n1425 VGND.n1342 146.25
R1296 VGND.n1425 VGND.n46 146.25
R1297 VGND.n1424 VGND.n1423 146.25
R1298 VGND.n1424 VGND.n47 146.25
R1299 VGND.n1422 VGND.n1344 146.25
R1300 VGND.n1344 VGND.n1343 146.25
R1301 VGND.n1421 VGND.n1420 146.25
R1302 VGND.n1420 VGND.n50 146.25
R1303 VGND.n1419 VGND.n1345 146.25
R1304 VGND.n1419 VGND.n51 146.25
R1305 VGND.n1418 VGND.n1417 146.25
R1306 VGND.n1418 VGND.n52 146.25
R1307 VGND.n1416 VGND.n1347 146.25
R1308 VGND.n1347 VGND.n1346 146.25
R1309 VGND.n1415 VGND.n1414 146.25
R1310 VGND.n1414 VGND.n55 146.25
R1311 VGND.n1413 VGND.n1348 146.25
R1312 VGND.n1413 VGND.n56 146.25
R1313 VGND.n1412 VGND.n1411 146.25
R1314 VGND.n1412 VGND.n57 146.25
R1315 VGND.n1410 VGND.n1350 146.25
R1316 VGND.n1350 VGND.n1349 146.25
R1317 VGND.n1409 VGND.n1408 146.25
R1318 VGND.n1408 VGND.n60 146.25
R1319 VGND.n1407 VGND.n1351 146.25
R1320 VGND.n1407 VGND.n61 146.25
R1321 VGND.n1406 VGND.n1405 146.25
R1322 VGND.n1406 VGND.n62 146.25
R1323 VGND.n1404 VGND.n1353 146.25
R1324 VGND.n1353 VGND.n1352 146.25
R1325 VGND.n1403 VGND.n1402 146.25
R1326 VGND.n1402 VGND.n65 146.25
R1327 VGND.n1401 VGND.n1354 146.25
R1328 VGND.n1401 VGND.n66 146.25
R1329 VGND.n1400 VGND.n1399 146.25
R1330 VGND.n1400 VGND.n67 146.25
R1331 VGND.n1398 VGND.n1356 146.25
R1332 VGND.n1356 VGND.n1355 146.25
R1333 VGND.n1397 VGND.n1396 146.25
R1334 VGND.n1396 VGND.n70 146.25
R1335 VGND.n1395 VGND.n1357 146.25
R1336 VGND.n1395 VGND.n71 146.25
R1337 VGND.n1394 VGND.n1393 146.25
R1338 VGND.n1394 VGND.n72 146.25
R1339 VGND.n1392 VGND.n1359 146.25
R1340 VGND.n1359 VGND.n1358 146.25
R1341 VGND.n1391 VGND.n1390 146.25
R1342 VGND.n1390 VGND.n75 146.25
R1343 VGND.n1389 VGND.n1360 146.25
R1344 VGND.n1389 VGND.n76 146.25
R1345 VGND.n1388 VGND.n1387 146.25
R1346 VGND.n1388 VGND.n77 146.25
R1347 VGND.n1386 VGND.n1362 146.25
R1348 VGND.n1362 VGND.n1361 146.25
R1349 VGND.n1385 VGND.n1384 146.25
R1350 VGND.n1384 VGND.n80 146.25
R1351 VGND.n1383 VGND.n1363 146.25
R1352 VGND.n1383 VGND.n81 146.25
R1353 VGND.n1382 VGND.n1381 146.25
R1354 VGND.n1382 VGND.n82 146.25
R1355 VGND.n1380 VGND.n1365 146.25
R1356 VGND.n1365 VGND.n1364 146.25
R1357 VGND.n1379 VGND.n1378 146.25
R1358 VGND.n1378 VGND.n85 146.25
R1359 VGND.n1377 VGND.n1366 146.25
R1360 VGND.n1377 VGND.n86 146.25
R1361 VGND.n1376 VGND.n1375 146.25
R1362 VGND.n1376 VGND.n87 146.25
R1363 VGND.n1374 VGND.n1368 146.25
R1364 VGND.n1368 VGND.n1367 146.25
R1365 VGND.n1373 VGND.n1372 146.25
R1366 VGND.n1372 VGND.n90 146.25
R1367 VGND.n1371 VGND.n1369 146.25
R1368 VGND.n1371 VGND.n91 146.25
R1369 VGND.n1370 VGND.n99 146.25
R1370 VGND.n1370 VGND.n92 146.25
R1371 VGND.n181 VGND.n98 146.25
R1372 VGND.n180 VGND.n94 146.25
R1373 VGND.n409 VGND.n184 146.25
R1374 VGND.n410 VGND.n179 146.25
R1375 VGND.n411 VGND.n187 146.25
R1376 VGND.n412 VGND.n178 146.25
R1377 VGND.n413 VGND.n190 146.25
R1378 VGND.n414 VGND.n177 146.25
R1379 VGND.n415 VGND.n193 146.25
R1380 VGND.n416 VGND.n176 146.25
R1381 VGND.n417 VGND.n196 146.25
R1382 VGND.n418 VGND.n175 146.25
R1383 VGND.n419 VGND.n199 146.25
R1384 VGND.n420 VGND.n174 146.25
R1385 VGND.n421 VGND.n202 146.25
R1386 VGND.n422 VGND.n173 146.25
R1387 VGND.n423 VGND.n205 146.25
R1388 VGND.n424 VGND.n172 146.25
R1389 VGND.n425 VGND.n208 146.25
R1390 VGND.n426 VGND.n171 146.25
R1391 VGND.n427 VGND.n211 146.25
R1392 VGND.n428 VGND.n170 146.25
R1393 VGND.n429 VGND.n214 146.25
R1394 VGND.n430 VGND.n169 146.25
R1395 VGND.n431 VGND.n217 146.25
R1396 VGND.n432 VGND.n168 146.25
R1397 VGND.n433 VGND.n220 146.25
R1398 VGND.n434 VGND.n167 146.25
R1399 VGND.n435 VGND.n223 146.25
R1400 VGND.n436 VGND.n166 146.25
R1401 VGND.n437 VGND.n226 146.25
R1402 VGND.n438 VGND.n165 146.25
R1403 VGND.n439 VGND.n229 146.25
R1404 VGND.n440 VGND.n164 146.25
R1405 VGND.n441 VGND.n232 146.25
R1406 VGND.n442 VGND.n163 146.25
R1407 VGND.n443 VGND.n235 146.25
R1408 VGND.n444 VGND.n162 146.25
R1409 VGND.n445 VGND.n238 146.25
R1410 VGND.n446 VGND.n161 146.25
R1411 VGND.n447 VGND.n241 146.25
R1412 VGND.n448 VGND.n160 146.25
R1413 VGND.n449 VGND.n244 146.25
R1414 VGND.n450 VGND.n159 146.25
R1415 VGND.n451 VGND.n247 146.25
R1416 VGND.n452 VGND.n158 146.25
R1417 VGND.n453 VGND.n250 146.25
R1418 VGND.n454 VGND.n157 146.25
R1419 VGND.n455 VGND.n253 146.25
R1420 VGND.n456 VGND.n156 146.25
R1421 VGND.n457 VGND.n256 146.25
R1422 VGND.n458 VGND.n155 146.25
R1423 VGND.n459 VGND.n259 146.25
R1424 VGND.n460 VGND.n154 146.25
R1425 VGND.n461 VGND.n262 146.25
R1426 VGND.n462 VGND.n153 146.25
R1427 VGND.n463 VGND.n265 146.25
R1428 VGND.n464 VGND.n152 146.25
R1429 VGND.n465 VGND.n268 146.25
R1430 VGND.n466 VGND.n151 146.25
R1431 VGND.n467 VGND.n271 146.25
R1432 VGND.n468 VGND.n150 146.25
R1433 VGND.n469 VGND.n274 146.25
R1434 VGND.n470 VGND.n149 146.25
R1435 VGND.n471 VGND.n277 146.25
R1436 VGND.n472 VGND.n148 146.25
R1437 VGND.n473 VGND.n280 146.25
R1438 VGND.n474 VGND.n147 146.25
R1439 VGND.n475 VGND.n283 146.25
R1440 VGND.n476 VGND.n146 146.25
R1441 VGND.n477 VGND.n286 146.25
R1442 VGND.n478 VGND.n145 146.25
R1443 VGND.n479 VGND.n289 146.25
R1444 VGND.n480 VGND.n144 146.25
R1445 VGND.n481 VGND.n292 146.25
R1446 VGND.n482 VGND.n143 146.25
R1447 VGND.n483 VGND.n295 146.25
R1448 VGND.n484 VGND.n142 146.25
R1449 VGND.n1485 VGND.n298 146.25
R1450 VGND.n1486 VGND.n141 146.25
R1451 VGND.n1487 VGND.n301 146.25
R1452 VGND.n1488 VGND.n140 146.25
R1453 VGND.n1489 VGND.n304 146.25
R1454 VGND.n1490 VGND.n139 146.25
R1455 VGND.n1491 VGND.n307 146.25
R1456 VGND.n1492 VGND.n138 146.25
R1457 VGND.n1493 VGND.n310 146.25
R1458 VGND.n1494 VGND.n137 146.25
R1459 VGND.n1495 VGND.n313 146.25
R1460 VGND.n1496 VGND.n136 146.25
R1461 VGND.n1497 VGND.n316 146.25
R1462 VGND.n1498 VGND.n135 146.25
R1463 VGND.n1499 VGND.n319 146.25
R1464 VGND.n1500 VGND.n134 146.25
R1465 VGND.n1501 VGND.n322 146.25
R1466 VGND.n1502 VGND.n133 146.25
R1467 VGND.n1503 VGND.n325 146.25
R1468 VGND.n1504 VGND.n132 146.25
R1469 VGND.n1505 VGND.n328 146.25
R1470 VGND.n1506 VGND.n131 146.25
R1471 VGND.n1507 VGND.n331 146.25
R1472 VGND.n1508 VGND.n130 146.25
R1473 VGND.n1509 VGND.n334 146.25
R1474 VGND.n1510 VGND.n129 146.25
R1475 VGND.n1511 VGND.n337 146.25
R1476 VGND.n1512 VGND.n128 146.25
R1477 VGND.n1513 VGND.n340 146.25
R1478 VGND.n1514 VGND.n127 146.25
R1479 VGND.n1515 VGND.n343 146.25
R1480 VGND.n1516 VGND.n126 146.25
R1481 VGND.n1517 VGND.n346 146.25
R1482 VGND.n1518 VGND.n125 146.25
R1483 VGND.n1519 VGND.n349 146.25
R1484 VGND.n1520 VGND.n124 146.25
R1485 VGND.n1521 VGND.n352 146.25
R1486 VGND.n1522 VGND.n123 146.25
R1487 VGND.n1523 VGND.n355 146.25
R1488 VGND.n1524 VGND.n122 146.25
R1489 VGND.n1525 VGND.n358 146.25
R1490 VGND.n1526 VGND.n121 146.25
R1491 VGND.n1527 VGND.n361 146.25
R1492 VGND.n1528 VGND.n120 146.25
R1493 VGND.n1529 VGND.n364 146.25
R1494 VGND.n1530 VGND.n119 146.25
R1495 VGND.n1531 VGND.n367 146.25
R1496 VGND.n1532 VGND.n118 146.25
R1497 VGND.n1533 VGND.n370 146.25
R1498 VGND.n1534 VGND.n117 146.25
R1499 VGND.n1535 VGND.n373 146.25
R1500 VGND.n1536 VGND.n116 146.25
R1501 VGND.n1537 VGND.n376 146.25
R1502 VGND.n1538 VGND.n115 146.25
R1503 VGND.n1539 VGND.n379 146.25
R1504 VGND.n1540 VGND.n114 146.25
R1505 VGND.n1541 VGND.n382 146.25
R1506 VGND.n1542 VGND.n113 146.25
R1507 VGND.n1543 VGND.n385 146.25
R1508 VGND.n1544 VGND.n112 146.25
R1509 VGND.n1545 VGND.n388 146.25
R1510 VGND.n1546 VGND.n111 146.25
R1511 VGND.n1547 VGND.n391 146.25
R1512 VGND.n1548 VGND.n110 146.25
R1513 VGND.n1549 VGND.n394 146.25
R1514 VGND.n1550 VGND.n109 146.25
R1515 VGND.n1551 VGND.n397 146.25
R1516 VGND.n1552 VGND.n108 146.25
R1517 VGND.n1553 VGND.n400 146.25
R1518 VGND.n1554 VGND.n107 146.25
R1519 VGND.n1555 VGND.n403 146.25
R1520 VGND.n1556 VGND.n106 146.25
R1521 VGND.n1557 VGND.n406 146.25
R1522 VGND.n1558 VGND.n105 146.25
R1523 VGND.n1560 VGND.n1559 146.25
R1524 VGND.n104 VGND.n100 146.25
R1525 VGND.n1563 VGND.n1562 146.25
R1526 VGND.n181 VGND.n95 146.25
R1527 VGND.n1570 VGND.n92 146.25
R1528 VGND.n1571 VGND.n91 146.25
R1529 VGND.n1572 VGND.n90 146.25
R1530 VGND.n1367 VGND.n88 146.25
R1531 VGND.n1576 VGND.n87 146.25
R1532 VGND.n1577 VGND.n86 146.25
R1533 VGND.n1578 VGND.n85 146.25
R1534 VGND.n1364 VGND.n83 146.25
R1535 VGND.n1582 VGND.n82 146.25
R1536 VGND.n1583 VGND.n81 146.25
R1537 VGND.n1584 VGND.n80 146.25
R1538 VGND.n1361 VGND.n78 146.25
R1539 VGND.n1588 VGND.n77 146.25
R1540 VGND.n1589 VGND.n76 146.25
R1541 VGND.n1590 VGND.n75 146.25
R1542 VGND.n1358 VGND.n73 146.25
R1543 VGND.n1594 VGND.n72 146.25
R1544 VGND.n1595 VGND.n71 146.25
R1545 VGND.n1596 VGND.n70 146.25
R1546 VGND.n1355 VGND.n68 146.25
R1547 VGND.n1600 VGND.n67 146.25
R1548 VGND.n1601 VGND.n66 146.25
R1549 VGND.n1602 VGND.n65 146.25
R1550 VGND.n1352 VGND.n63 146.25
R1551 VGND.n1606 VGND.n62 146.25
R1552 VGND.n1607 VGND.n61 146.25
R1553 VGND.n1608 VGND.n60 146.25
R1554 VGND.n1349 VGND.n58 146.25
R1555 VGND.n1612 VGND.n57 146.25
R1556 VGND.n1613 VGND.n56 146.25
R1557 VGND.n1614 VGND.n55 146.25
R1558 VGND.n1346 VGND.n53 146.25
R1559 VGND.n1618 VGND.n52 146.25
R1560 VGND.n1619 VGND.n51 146.25
R1561 VGND.n1620 VGND.n50 146.25
R1562 VGND.n1343 VGND.n48 146.25
R1563 VGND.n1624 VGND.n47 146.25
R1564 VGND.n1625 VGND.n46 146.25
R1565 VGND.n1626 VGND.n45 146.25
R1566 VGND.n1340 VGND.n43 146.25
R1567 VGND.n1630 VGND.n42 146.25
R1568 VGND.n1631 VGND.n41 146.25
R1569 VGND.n1632 VGND.n40 146.25
R1570 VGND.n1337 VGND.n38 146.25
R1571 VGND.n1636 VGND.n37 146.25
R1572 VGND.n1637 VGND.n36 146.25
R1573 VGND.n1638 VGND.n35 146.25
R1574 VGND.n1334 VGND.n33 146.25
R1575 VGND.n1642 VGND.n32 146.25
R1576 VGND.n1643 VGND.n31 146.25
R1577 VGND.n1644 VGND.n30 146.25
R1578 VGND.n1331 VGND.n28 146.25
R1579 VGND.n1648 VGND.n27 146.25
R1580 VGND.n1649 VGND.n26 146.25
R1581 VGND.n1650 VGND.n25 146.25
R1582 VGND.n1328 VGND.n23 146.25
R1583 VGND.n1654 VGND.n22 146.25
R1584 VGND.n1655 VGND.n21 146.25
R1585 VGND.n1656 VGND.n20 146.25
R1586 VGND.n1325 VGND.n18 146.25
R1587 VGND.n1660 VGND.n17 146.25
R1588 VGND.n1661 VGND.n16 146.25
R1589 VGND.n1662 VGND.n15 146.25
R1590 VGND.n1322 VGND.n13 146.25
R1591 VGND.n1666 VGND.n12 146.25
R1592 VGND.n1667 VGND.n11 146.25
R1593 VGND.n1668 VGND.n10 146.25
R1594 VGND.n1319 VGND.n8 146.25
R1595 VGND.n1672 VGND.n7 146.25
R1596 VGND.n1673 VGND.n6 146.25
R1597 VGND.n1674 VGND.n5 146.25
R1598 VGND.n1316 VGND.n1315 146.25
R1599 VGND.n1314 VGND.n488 146.25
R1600 VGND.n493 VGND.n489 146.25
R1601 VGND.n1310 VGND.n1309 146.25
R1602 VGND.n492 VGND.n491 146.25
R1603 VGND.n1300 VGND.n1299 146.25
R1604 VGND.n499 VGND.n498 146.25
R1605 VGND.n1295 VGND.n1294 146.25
R1606 VGND.n502 VGND.n501 146.25
R1607 VGND.n1288 VGND.n1287 146.25
R1608 VGND.n510 VGND.n506 146.25
R1609 VGND.n1283 VGND.n1282 146.25
R1610 VGND.n509 VGND.n508 146.25
R1611 VGND.n1276 VGND.n1275 146.25
R1612 VGND.n515 VGND.n514 146.25
R1613 VGND.n1271 VGND.n1270 146.25
R1614 VGND.n518 VGND.n517 146.25
R1615 VGND.n1264 VGND.n1263 146.25
R1616 VGND.n523 VGND.n522 146.25
R1617 VGND.n1259 VGND.n1258 146.25
R1618 VGND.n530 VGND.n525 146.25
R1619 VGND.n1252 VGND.n1251 146.25
R1620 VGND.n531 VGND.n529 146.25
R1621 VGND.n1247 VGND.n1246 146.25
R1622 VGND.n534 VGND.n533 146.25
R1623 VGND.n1240 VGND.n1239 146.25
R1624 VGND.n539 VGND.n538 146.25
R1625 VGND.n1235 VGND.n1234 146.25
R1626 VGND.n542 VGND.n541 146.25
R1627 VGND.n1228 VGND.n1227 146.25
R1628 VGND.n550 VGND.n546 146.25
R1629 VGND.n1223 VGND.n1222 146.25
R1630 VGND.n549 VGND.n548 146.25
R1631 VGND.n1216 VGND.n1215 146.25
R1632 VGND.n555 VGND.n554 146.25
R1633 VGND.n1211 VGND.n1210 146.25
R1634 VGND.n558 VGND.n557 146.25
R1635 VGND.n1204 VGND.n1203 146.25
R1636 VGND.n563 VGND.n562 146.25
R1637 VGND.n1199 VGND.n1198 146.25
R1638 VGND.n570 VGND.n565 146.25
R1639 VGND.n1192 VGND.n1191 146.25
R1640 VGND.n571 VGND.n569 146.25
R1641 VGND.n1187 VGND.n1186 146.25
R1642 VGND.n574 VGND.n573 146.25
R1643 VGND.n1180 VGND.n1179 146.25
R1644 VGND.n579 VGND.n578 146.25
R1645 VGND.n1175 VGND.n1174 146.25
R1646 VGND.n582 VGND.n581 146.25
R1647 VGND.n1168 VGND.n1167 146.25
R1648 VGND.n590 VGND.n586 146.25
R1649 VGND.n1163 VGND.n1162 146.25
R1650 VGND.n589 VGND.n588 146.25
R1651 VGND.n1156 VGND.n1155 146.25
R1652 VGND.n595 VGND.n594 146.25
R1653 VGND.n1151 VGND.n1150 146.25
R1654 VGND.n598 VGND.n597 146.25
R1655 VGND.n1144 VGND.n1143 146.25
R1656 VGND.n603 VGND.n602 146.25
R1657 VGND.n1139 VGND.n1138 146.25
R1658 VGND.n610 VGND.n605 146.25
R1659 VGND.n1132 VGND.n1131 146.25
R1660 VGND.n611 VGND.n609 146.25
R1661 VGND.n1127 VGND.n1126 146.25
R1662 VGND.n614 VGND.n613 146.25
R1663 VGND.n1120 VGND.n1119 146.25
R1664 VGND.n619 VGND.n618 146.25
R1665 VGND.n1115 VGND.n1114 146.25
R1666 VGND.n622 VGND.n621 146.25
R1667 VGND.n1108 VGND.n1107 146.25
R1668 VGND.n937 VGND.n627 146.25
R1669 VGND.n1102 VGND.n630 146.25
R1670 VGND.t15 VGND.n3 146.25
R1671 VGND.n1570 VGND.n1569 146.25
R1672 VGND.n1571 VGND.n89 146.25
R1673 VGND.n1573 VGND.n1572 146.25
R1674 VGND.n1574 VGND.n88 146.25
R1675 VGND.n1576 VGND.n1575 146.25
R1676 VGND.n1577 VGND.n84 146.25
R1677 VGND.n1579 VGND.n1578 146.25
R1678 VGND.n1580 VGND.n83 146.25
R1679 VGND.n1582 VGND.n1581 146.25
R1680 VGND.n1583 VGND.n79 146.25
R1681 VGND.n1585 VGND.n1584 146.25
R1682 VGND.n1586 VGND.n78 146.25
R1683 VGND.n1588 VGND.n1587 146.25
R1684 VGND.n1589 VGND.n74 146.25
R1685 VGND.n1591 VGND.n1590 146.25
R1686 VGND.n1592 VGND.n73 146.25
R1687 VGND.n1594 VGND.n1593 146.25
R1688 VGND.n1595 VGND.n69 146.25
R1689 VGND.n1597 VGND.n1596 146.25
R1690 VGND.n1598 VGND.n68 146.25
R1691 VGND.n1600 VGND.n1599 146.25
R1692 VGND.n1601 VGND.n64 146.25
R1693 VGND.n1603 VGND.n1602 146.25
R1694 VGND.n1604 VGND.n63 146.25
R1695 VGND.n1606 VGND.n1605 146.25
R1696 VGND.n1607 VGND.n59 146.25
R1697 VGND.n1609 VGND.n1608 146.25
R1698 VGND.n1610 VGND.n58 146.25
R1699 VGND.n1612 VGND.n1611 146.25
R1700 VGND.n1613 VGND.n54 146.25
R1701 VGND.n1615 VGND.n1614 146.25
R1702 VGND.n1616 VGND.n53 146.25
R1703 VGND.n1618 VGND.n1617 146.25
R1704 VGND.n1619 VGND.n49 146.25
R1705 VGND.n1621 VGND.n1620 146.25
R1706 VGND.n1622 VGND.n48 146.25
R1707 VGND.n1624 VGND.n1623 146.25
R1708 VGND.n1625 VGND.n44 146.25
R1709 VGND.n1627 VGND.n1626 146.25
R1710 VGND.n1628 VGND.n43 146.25
R1711 VGND.n1630 VGND.n1629 146.25
R1712 VGND.n1631 VGND.n39 146.25
R1713 VGND.n1633 VGND.n1632 146.25
R1714 VGND.n1634 VGND.n38 146.25
R1715 VGND.n1636 VGND.n1635 146.25
R1716 VGND.n1637 VGND.n34 146.25
R1717 VGND.n1639 VGND.n1638 146.25
R1718 VGND.n1640 VGND.n33 146.25
R1719 VGND.n1642 VGND.n1641 146.25
R1720 VGND.n1643 VGND.n29 146.25
R1721 VGND.n1645 VGND.n1644 146.25
R1722 VGND.n1646 VGND.n28 146.25
R1723 VGND.n1648 VGND.n1647 146.25
R1724 VGND.n1649 VGND.n24 146.25
R1725 VGND.n1651 VGND.n1650 146.25
R1726 VGND.n1652 VGND.n23 146.25
R1727 VGND.n1654 VGND.n1653 146.25
R1728 VGND.n1655 VGND.n19 146.25
R1729 VGND.n1657 VGND.n1656 146.25
R1730 VGND.n1658 VGND.n18 146.25
R1731 VGND.n1660 VGND.n1659 146.25
R1732 VGND.n1661 VGND.n14 146.25
R1733 VGND.n1663 VGND.n1662 146.25
R1734 VGND.n1664 VGND.n13 146.25
R1735 VGND.n1666 VGND.n1665 146.25
R1736 VGND.n1667 VGND.n9 146.25
R1737 VGND.n1669 VGND.n1668 146.25
R1738 VGND.n1670 VGND.n8 146.25
R1739 VGND.n1672 VGND.n1671 146.25
R1740 VGND.n1673 VGND.n4 146.25
R1741 VGND.n1675 VGND.n1674 146.25
R1742 VGND.n1676 VGND.n3 146.25
R1743 VGND.n1315 VGND.n2 146.25
R1744 VGND.n1314 VGND.n1313 146.25
R1745 VGND.n1312 VGND.n489 146.25
R1746 VGND.n1311 VGND.n1310 146.25
R1747 VGND.n491 VGND.n490 146.25
R1748 VGND.n1299 VGND.n1298 146.25
R1749 VGND.n1297 VGND.n499 146.25
R1750 VGND.n1296 VGND.n1295 146.25
R1751 VGND.n501 VGND.n500 146.25
R1752 VGND.n1287 VGND.n1286 146.25
R1753 VGND.n1285 VGND.n506 146.25
R1754 VGND.n1284 VGND.n1283 146.25
R1755 VGND.n508 VGND.n507 146.25
R1756 VGND.n1275 VGND.n1274 146.25
R1757 VGND.n1273 VGND.n515 146.25
R1758 VGND.n1272 VGND.n1271 146.25
R1759 VGND.n517 VGND.n516 146.25
R1760 VGND.n1263 VGND.n1262 146.25
R1761 VGND.n1261 VGND.n523 146.25
R1762 VGND.n1260 VGND.n1259 146.25
R1763 VGND.n525 VGND.n524 146.25
R1764 VGND.n1251 VGND.n1250 146.25
R1765 VGND.n1249 VGND.n531 146.25
R1766 VGND.n1248 VGND.n1247 146.25
R1767 VGND.n533 VGND.n532 146.25
R1768 VGND.n1239 VGND.n1238 146.25
R1769 VGND.n1237 VGND.n539 146.25
R1770 VGND.n1236 VGND.n1235 146.25
R1771 VGND.n541 VGND.n540 146.25
R1772 VGND.n1227 VGND.n1226 146.25
R1773 VGND.n1225 VGND.n546 146.25
R1774 VGND.n1224 VGND.n1223 146.25
R1775 VGND.n548 VGND.n547 146.25
R1776 VGND.n1215 VGND.n1214 146.25
R1777 VGND.n1213 VGND.n555 146.25
R1778 VGND.n1212 VGND.n1211 146.25
R1779 VGND.n557 VGND.n556 146.25
R1780 VGND.n1203 VGND.n1202 146.25
R1781 VGND.n1201 VGND.n563 146.25
R1782 VGND.n1200 VGND.n1199 146.25
R1783 VGND.n565 VGND.n564 146.25
R1784 VGND.n1191 VGND.n1190 146.25
R1785 VGND.n1189 VGND.n571 146.25
R1786 VGND.n1188 VGND.n1187 146.25
R1787 VGND.n573 VGND.n572 146.25
R1788 VGND.n1179 VGND.n1178 146.25
R1789 VGND.n1177 VGND.n579 146.25
R1790 VGND.n1176 VGND.n1175 146.25
R1791 VGND.n581 VGND.n580 146.25
R1792 VGND.n1167 VGND.n1166 146.25
R1793 VGND.n1165 VGND.n586 146.25
R1794 VGND.n1164 VGND.n1163 146.25
R1795 VGND.n588 VGND.n587 146.25
R1796 VGND.n1155 VGND.n1154 146.25
R1797 VGND.n1153 VGND.n595 146.25
R1798 VGND.n1152 VGND.n1151 146.25
R1799 VGND.n597 VGND.n596 146.25
R1800 VGND.n1143 VGND.n1142 146.25
R1801 VGND.n1141 VGND.n603 146.25
R1802 VGND.n1140 VGND.n1139 146.25
R1803 VGND.n605 VGND.n604 146.25
R1804 VGND.n1131 VGND.n1130 146.25
R1805 VGND.n1129 VGND.n611 146.25
R1806 VGND.n1128 VGND.n1127 146.25
R1807 VGND.n613 VGND.n612 146.25
R1808 VGND.n1119 VGND.n1118 146.25
R1809 VGND.n1117 VGND.n619 146.25
R1810 VGND.n1116 VGND.n1115 146.25
R1811 VGND.n621 VGND.n620 146.25
R1812 VGND.n1107 VGND.n1106 146.25
R1813 VGND.n1105 VGND.n627 146.25
R1814 VGND.n942 VGND.n941 65.1484
R1815 VGND.n1568 VGND.n1567 65.1484
R1816 VGND.n1565 VGND.n1564 65.1478
R1817 VGND.n1104 VGND.n1103 65.1478
R1818 VGND.n1562 VGND.n101 60.4138
R1819 VGND.n180 VGND.n93 60.4138
R1820 VGND.n1098 VGND.n861 60.4138
R1821 VGND.n1101 VGND.n1100 60.4138
R1822 VGND.n1109 VGND.n625 47.2805
R1823 VGND.n1109 VGND.n623 47.2805
R1824 VGND.n1113 VGND.n623 47.2805
R1825 VGND.n1113 VGND.n617 47.2805
R1826 VGND.n1121 VGND.n617 47.2805
R1827 VGND.n1121 VGND.n615 47.2805
R1828 VGND.n1125 VGND.n615 47.2805
R1829 VGND.n1125 VGND.n608 47.2805
R1830 VGND.n1133 VGND.n608 47.2805
R1831 VGND.n1133 VGND.n606 47.2805
R1832 VGND.n1137 VGND.n606 47.2805
R1833 VGND.n1137 VGND.n601 47.2805
R1834 VGND.n1145 VGND.n601 47.2805
R1835 VGND.n1145 VGND.n599 47.2805
R1836 VGND.n1149 VGND.n599 47.2805
R1837 VGND.n1149 VGND.n593 47.2805
R1838 VGND.n1157 VGND.n593 47.2805
R1839 VGND.n1157 VGND.n591 47.2805
R1840 VGND.n1161 VGND.n591 47.2805
R1841 VGND.n1161 VGND.n585 47.2805
R1842 VGND.n1169 VGND.n585 47.2805
R1843 VGND.n1169 VGND.n583 47.2805
R1844 VGND.n1173 VGND.n583 47.2805
R1845 VGND.n1173 VGND.n577 47.2805
R1846 VGND.n1181 VGND.n577 47.2805
R1847 VGND.n1181 VGND.n575 47.2805
R1848 VGND.n1185 VGND.n575 47.2805
R1849 VGND.n1185 VGND.n568 47.2805
R1850 VGND.n1193 VGND.n568 47.2805
R1851 VGND.n1193 VGND.n566 47.2805
R1852 VGND.n1197 VGND.n566 47.2805
R1853 VGND.n1197 VGND.n561 47.2805
R1854 VGND.n1205 VGND.n561 47.2805
R1855 VGND.n1205 VGND.n559 47.2805
R1856 VGND.n1209 VGND.n559 47.2805
R1857 VGND.n1209 VGND.n553 47.2805
R1858 VGND.n1217 VGND.n553 47.2805
R1859 VGND.n1217 VGND.n551 47.2805
R1860 VGND.n1221 VGND.n551 47.2805
R1861 VGND.n1221 VGND.n545 47.2805
R1862 VGND.n1229 VGND.n545 47.2805
R1863 VGND.n1229 VGND.n543 47.2805
R1864 VGND.n1233 VGND.n543 47.2805
R1865 VGND.n1233 VGND.n537 47.2805
R1866 VGND.n1241 VGND.n537 47.2805
R1867 VGND.n1241 VGND.n535 47.2805
R1868 VGND.n1245 VGND.n535 47.2805
R1869 VGND.n1245 VGND.n528 47.2805
R1870 VGND.n1253 VGND.n528 47.2805
R1871 VGND.n1253 VGND.n526 47.2805
R1872 VGND.n1257 VGND.n526 47.2805
R1873 VGND.n1257 VGND.n521 47.2805
R1874 VGND.n1265 VGND.n521 47.2805
R1875 VGND.n1265 VGND.n519 47.2805
R1876 VGND.n1269 VGND.n519 47.2805
R1877 VGND.n1269 VGND.n513 47.2805
R1878 VGND.n1277 VGND.n513 47.2805
R1879 VGND.n1277 VGND.n511 47.2805
R1880 VGND.n1281 VGND.n511 47.2805
R1881 VGND.n1281 VGND.n505 47.2805
R1882 VGND.n1289 VGND.n505 47.2805
R1883 VGND.n1289 VGND.n503 47.2805
R1884 VGND.n1293 VGND.n503 47.2805
R1885 VGND.n1293 VGND.n497 47.2805
R1886 VGND.n1301 VGND.n497 47.2805
R1887 VGND.n1301 VGND.n494 47.2805
R1888 VGND.n1308 VGND.n494 47.2805
R1889 VGND.n1308 VGND.n495 47.2805
R1890 VGND.n1304 VGND.n495 47.2805
R1891 VGND.n1304 VGND.n487 47.2805
R1892 VGND.n1317 VGND.n487 47.2805
R1893 VGND.n1474 VGND.n1317 47.2805
R1894 VGND.n1474 VGND.n1473 47.2805
R1895 VGND.n1473 VGND.n1472 47.2805
R1896 VGND.n1472 VGND.n1320 47.2805
R1897 VGND.n1468 VGND.n1320 47.2805
R1898 VGND.n1468 VGND.n1467 47.2805
R1899 VGND.n1467 VGND.n1466 47.2805
R1900 VGND.n1466 VGND.n1323 47.2805
R1901 VGND.n1462 VGND.n1323 47.2805
R1902 VGND.n1462 VGND.n1461 47.2805
R1903 VGND.n1461 VGND.n1460 47.2805
R1904 VGND.n1460 VGND.n1326 47.2805
R1905 VGND.n1456 VGND.n1326 47.2805
R1906 VGND.n1456 VGND.n1455 47.2805
R1907 VGND.n1455 VGND.n1454 47.2805
R1908 VGND.n1454 VGND.n1329 47.2805
R1909 VGND.n1450 VGND.n1329 47.2805
R1910 VGND.n1450 VGND.n1449 47.2805
R1911 VGND.n1449 VGND.n1448 47.2805
R1912 VGND.n1448 VGND.n1332 47.2805
R1913 VGND.n1444 VGND.n1332 47.2805
R1914 VGND.n1444 VGND.n1443 47.2805
R1915 VGND.n1443 VGND.n1442 47.2805
R1916 VGND.n1442 VGND.n1335 47.2805
R1917 VGND.n1438 VGND.n1335 47.2805
R1918 VGND.n1438 VGND.n1437 47.2805
R1919 VGND.n1437 VGND.n1436 47.2805
R1920 VGND.n1436 VGND.n1338 47.2805
R1921 VGND.n1432 VGND.n1338 47.2805
R1922 VGND.n1432 VGND.n1431 47.2805
R1923 VGND.n1431 VGND.n1430 47.2805
R1924 VGND.n1430 VGND.n1341 47.2805
R1925 VGND.n1426 VGND.n1341 47.2805
R1926 VGND.n1426 VGND.n1425 47.2805
R1927 VGND.n1425 VGND.n1424 47.2805
R1928 VGND.n1424 VGND.n1344 47.2805
R1929 VGND.n1420 VGND.n1344 47.2805
R1930 VGND.n1420 VGND.n1419 47.2805
R1931 VGND.n1419 VGND.n1418 47.2805
R1932 VGND.n1418 VGND.n1347 47.2805
R1933 VGND.n1414 VGND.n1347 47.2805
R1934 VGND.n1414 VGND.n1413 47.2805
R1935 VGND.n1413 VGND.n1412 47.2805
R1936 VGND.n1412 VGND.n1350 47.2805
R1937 VGND.n1408 VGND.n1350 47.2805
R1938 VGND.n1408 VGND.n1407 47.2805
R1939 VGND.n1407 VGND.n1406 47.2805
R1940 VGND.n1406 VGND.n1353 47.2805
R1941 VGND.n1402 VGND.n1353 47.2805
R1942 VGND.n1402 VGND.n1401 47.2805
R1943 VGND.n1401 VGND.n1400 47.2805
R1944 VGND.n1400 VGND.n1356 47.2805
R1945 VGND.n1396 VGND.n1356 47.2805
R1946 VGND.n1396 VGND.n1395 47.2805
R1947 VGND.n1395 VGND.n1394 47.2805
R1948 VGND.n1394 VGND.n1359 47.2805
R1949 VGND.n1390 VGND.n1359 47.2805
R1950 VGND.n1390 VGND.n1389 47.2805
R1951 VGND.n1389 VGND.n1388 47.2805
R1952 VGND.n1388 VGND.n1362 47.2805
R1953 VGND.n1384 VGND.n1362 47.2805
R1954 VGND.n1384 VGND.n1383 47.2805
R1955 VGND.n1383 VGND.n1382 47.2805
R1956 VGND.n1382 VGND.n1365 47.2805
R1957 VGND.n1378 VGND.n1365 47.2805
R1958 VGND.n1378 VGND.n1377 47.2805
R1959 VGND.n1377 VGND.n1376 47.2805
R1960 VGND.n1376 VGND.n1368 47.2805
R1961 VGND.n1372 VGND.n1368 47.2805
R1962 VGND.n1372 VGND.n1371 47.2805
R1963 VGND.n1371 VGND.n1370 47.2805
R1964 VGND.n1107 VGND.n627 47.2805
R1965 VGND.n1107 VGND.n621 47.2805
R1966 VGND.n1115 VGND.n621 47.2805
R1967 VGND.n1115 VGND.n619 47.2805
R1968 VGND.n1119 VGND.n619 47.2805
R1969 VGND.n1119 VGND.n613 47.2805
R1970 VGND.n1127 VGND.n613 47.2805
R1971 VGND.n1127 VGND.n611 47.2805
R1972 VGND.n1131 VGND.n611 47.2805
R1973 VGND.n1131 VGND.n605 47.2805
R1974 VGND.n1139 VGND.n605 47.2805
R1975 VGND.n1139 VGND.n603 47.2805
R1976 VGND.n1143 VGND.n603 47.2805
R1977 VGND.n1143 VGND.n597 47.2805
R1978 VGND.n1151 VGND.n597 47.2805
R1979 VGND.n1151 VGND.n595 47.2805
R1980 VGND.n1155 VGND.n595 47.2805
R1981 VGND.n1155 VGND.n588 47.2805
R1982 VGND.n1163 VGND.n588 47.2805
R1983 VGND.n1163 VGND.n586 47.2805
R1984 VGND.n1167 VGND.n586 47.2805
R1985 VGND.n1167 VGND.n581 47.2805
R1986 VGND.n1175 VGND.n581 47.2805
R1987 VGND.n1175 VGND.n579 47.2805
R1988 VGND.n1179 VGND.n579 47.2805
R1989 VGND.n1179 VGND.n573 47.2805
R1990 VGND.n1187 VGND.n573 47.2805
R1991 VGND.n1187 VGND.n571 47.2805
R1992 VGND.n1191 VGND.n571 47.2805
R1993 VGND.n1191 VGND.n565 47.2805
R1994 VGND.n1199 VGND.n565 47.2805
R1995 VGND.n1199 VGND.n563 47.2805
R1996 VGND.n1203 VGND.n563 47.2805
R1997 VGND.n1203 VGND.n557 47.2805
R1998 VGND.n1211 VGND.n557 47.2805
R1999 VGND.n1211 VGND.n555 47.2805
R2000 VGND.n1215 VGND.n555 47.2805
R2001 VGND.n1215 VGND.n548 47.2805
R2002 VGND.n1223 VGND.n548 47.2805
R2003 VGND.n1223 VGND.n546 47.2805
R2004 VGND.n1227 VGND.n546 47.2805
R2005 VGND.n1227 VGND.n541 47.2805
R2006 VGND.n1235 VGND.n541 47.2805
R2007 VGND.n1235 VGND.n539 47.2805
R2008 VGND.n1239 VGND.n539 47.2805
R2009 VGND.n1239 VGND.n533 47.2805
R2010 VGND.n1247 VGND.n533 47.2805
R2011 VGND.n1247 VGND.n531 47.2805
R2012 VGND.n1251 VGND.n531 47.2805
R2013 VGND.n1251 VGND.n525 47.2805
R2014 VGND.n1259 VGND.n525 47.2805
R2015 VGND.n1259 VGND.n523 47.2805
R2016 VGND.n1263 VGND.n523 47.2805
R2017 VGND.n1263 VGND.n517 47.2805
R2018 VGND.n1271 VGND.n517 47.2805
R2019 VGND.n1271 VGND.n515 47.2805
R2020 VGND.n1275 VGND.n515 47.2805
R2021 VGND.n1275 VGND.n508 47.2805
R2022 VGND.n1283 VGND.n508 47.2805
R2023 VGND.n1283 VGND.n506 47.2805
R2024 VGND.n1287 VGND.n506 47.2805
R2025 VGND.n1287 VGND.n501 47.2805
R2026 VGND.n1295 VGND.n501 47.2805
R2027 VGND.n1295 VGND.n499 47.2805
R2028 VGND.n1299 VGND.n499 47.2805
R2029 VGND.n1299 VGND.n491 47.2805
R2030 VGND.n1310 VGND.n491 47.2805
R2031 VGND.n1310 VGND.n489 47.2805
R2032 VGND.n1314 VGND.n489 47.2805
R2033 VGND.n1315 VGND.n1314 47.2805
R2034 VGND.n1315 VGND.n3 47.2805
R2035 VGND.n1674 VGND.n3 47.2805
R2036 VGND.n1674 VGND.n1673 47.2805
R2037 VGND.n1673 VGND.n1672 47.2805
R2038 VGND.n1672 VGND.n8 47.2805
R2039 VGND.n1668 VGND.n8 47.2805
R2040 VGND.n1668 VGND.n1667 47.2805
R2041 VGND.n1667 VGND.n1666 47.2805
R2042 VGND.n1666 VGND.n13 47.2805
R2043 VGND.n1662 VGND.n13 47.2805
R2044 VGND.n1662 VGND.n1661 47.2805
R2045 VGND.n1661 VGND.n1660 47.2805
R2046 VGND.n1660 VGND.n18 47.2805
R2047 VGND.n1656 VGND.n18 47.2805
R2048 VGND.n1656 VGND.n1655 47.2805
R2049 VGND.n1655 VGND.n1654 47.2805
R2050 VGND.n1654 VGND.n23 47.2805
R2051 VGND.n1650 VGND.n23 47.2805
R2052 VGND.n1650 VGND.n1649 47.2805
R2053 VGND.n1649 VGND.n1648 47.2805
R2054 VGND.n1648 VGND.n28 47.2805
R2055 VGND.n1644 VGND.n28 47.2805
R2056 VGND.n1644 VGND.n1643 47.2805
R2057 VGND.n1643 VGND.n1642 47.2805
R2058 VGND.n1642 VGND.n33 47.2805
R2059 VGND.n1638 VGND.n33 47.2805
R2060 VGND.n1638 VGND.n1637 47.2805
R2061 VGND.n1637 VGND.n1636 47.2805
R2062 VGND.n1636 VGND.n38 47.2805
R2063 VGND.n1632 VGND.n38 47.2805
R2064 VGND.n1632 VGND.n1631 47.2805
R2065 VGND.n1631 VGND.n1630 47.2805
R2066 VGND.n1630 VGND.n43 47.2805
R2067 VGND.n1626 VGND.n43 47.2805
R2068 VGND.n1626 VGND.n1625 47.2805
R2069 VGND.n1625 VGND.n1624 47.2805
R2070 VGND.n1624 VGND.n48 47.2805
R2071 VGND.n1620 VGND.n48 47.2805
R2072 VGND.n1620 VGND.n1619 47.2805
R2073 VGND.n1619 VGND.n1618 47.2805
R2074 VGND.n1618 VGND.n53 47.2805
R2075 VGND.n1614 VGND.n53 47.2805
R2076 VGND.n1614 VGND.n1613 47.2805
R2077 VGND.n1613 VGND.n1612 47.2805
R2078 VGND.n1612 VGND.n58 47.2805
R2079 VGND.n1608 VGND.n58 47.2805
R2080 VGND.n1608 VGND.n1607 47.2805
R2081 VGND.n1607 VGND.n1606 47.2805
R2082 VGND.n1606 VGND.n63 47.2805
R2083 VGND.n1602 VGND.n63 47.2805
R2084 VGND.n1602 VGND.n1601 47.2805
R2085 VGND.n1601 VGND.n1600 47.2805
R2086 VGND.n1600 VGND.n68 47.2805
R2087 VGND.n1596 VGND.n68 47.2805
R2088 VGND.n1596 VGND.n1595 47.2805
R2089 VGND.n1595 VGND.n1594 47.2805
R2090 VGND.n1594 VGND.n73 47.2805
R2091 VGND.n1590 VGND.n73 47.2805
R2092 VGND.n1590 VGND.n1589 47.2805
R2093 VGND.n1589 VGND.n1588 47.2805
R2094 VGND.n1588 VGND.n78 47.2805
R2095 VGND.n1584 VGND.n78 47.2805
R2096 VGND.n1584 VGND.n1583 47.2805
R2097 VGND.n1583 VGND.n1582 47.2805
R2098 VGND.n1582 VGND.n83 47.2805
R2099 VGND.n1578 VGND.n83 47.2805
R2100 VGND.n1578 VGND.n1577 47.2805
R2101 VGND.n1577 VGND.n1576 47.2805
R2102 VGND.n1576 VGND.n88 47.2805
R2103 VGND.n1572 VGND.n88 47.2805
R2104 VGND.n1572 VGND.n1571 47.2805
R2105 VGND.n1571 VGND.n1570 47.2805
R2106 VGND.n1108 VGND.n622 26.7302
R2107 VGND.n1114 VGND.n622 26.7302
R2108 VGND.n1114 VGND.n618 26.7302
R2109 VGND.n1120 VGND.n618 26.7302
R2110 VGND.n1126 VGND.n614 26.7302
R2111 VGND.n1126 VGND.n609 26.7302
R2112 VGND.n1132 VGND.n609 26.7302
R2113 VGND.n1132 VGND.n610 26.7302
R2114 VGND.n1138 VGND.n602 26.7302
R2115 VGND.n1144 VGND.n602 26.7302
R2116 VGND.n1144 VGND.n598 26.7302
R2117 VGND.n1150 VGND.n598 26.7302
R2118 VGND.n1156 VGND.n594 26.7302
R2119 VGND.n1156 VGND.n589 26.7302
R2120 VGND.n1162 VGND.n589 26.7302
R2121 VGND.n1162 VGND.n590 26.7302
R2122 VGND.n1168 VGND.n582 26.7302
R2123 VGND.n1174 VGND.n582 26.7302
R2124 VGND.n1174 VGND.n578 26.7302
R2125 VGND.n1180 VGND.n578 26.7302
R2126 VGND.n1186 VGND.n574 26.7302
R2127 VGND.n1186 VGND.n569 26.7302
R2128 VGND.n1192 VGND.n569 26.7302
R2129 VGND.n1192 VGND.n570 26.7302
R2130 VGND.n1198 VGND.n562 26.7302
R2131 VGND.n1204 VGND.n562 26.7302
R2132 VGND.n1204 VGND.n558 26.7302
R2133 VGND.n1210 VGND.n558 26.7302
R2134 VGND.n1216 VGND.n554 26.7302
R2135 VGND.n1216 VGND.n549 26.7302
R2136 VGND.n1222 VGND.n549 26.7302
R2137 VGND.n1222 VGND.n550 26.7302
R2138 VGND.n1228 VGND.n542 26.7302
R2139 VGND.n1234 VGND.n542 26.7302
R2140 VGND.n1234 VGND.n538 26.7302
R2141 VGND.n1240 VGND.n538 26.7302
R2142 VGND.n1246 VGND.n534 26.7302
R2143 VGND.n1246 VGND.n529 26.7302
R2144 VGND.n1252 VGND.n529 26.7302
R2145 VGND.n1252 VGND.n530 26.7302
R2146 VGND.n1258 VGND.n522 26.7302
R2147 VGND.n1264 VGND.n522 26.7302
R2148 VGND.n1264 VGND.n518 26.7302
R2149 VGND.n1270 VGND.n518 26.7302
R2150 VGND.n1276 VGND.n514 26.7302
R2151 VGND.n1276 VGND.n509 26.7302
R2152 VGND.n1282 VGND.n509 26.7302
R2153 VGND.n1282 VGND.n510 26.7302
R2154 VGND.n1288 VGND.n502 26.7302
R2155 VGND.n1294 VGND.n502 26.7302
R2156 VGND.n1294 VGND.n498 26.7302
R2157 VGND.n1300 VGND.n498 26.7302
R2158 VGND.n1309 VGND.n492 26.7302
R2159 VGND.n1309 VGND.n493 26.7302
R2160 VGND.n493 VGND.n488 26.7302
R2161 VGND.n1316 VGND.n488 26.7302
R2162 VGND.t15 VGND.n1316 26.7302
R2163 VGND.t15 VGND.n5 26.7302
R2164 VGND.n6 VGND.n5 26.7302
R2165 VGND.n7 VGND.n6 26.7302
R2166 VGND.n1319 VGND.n7 26.7302
R2167 VGND.n1319 VGND.n10 26.7302
R2168 VGND.n12 VGND.n11 26.7302
R2169 VGND.n1322 VGND.n12 26.7302
R2170 VGND.n1322 VGND.n15 26.7302
R2171 VGND.n16 VGND.n15 26.7302
R2172 VGND.n1325 VGND.n17 26.7302
R2173 VGND.n1325 VGND.n20 26.7302
R2174 VGND.n21 VGND.n20 26.7302
R2175 VGND.n22 VGND.n21 26.7302
R2176 VGND.n1328 VGND.n25 26.7302
R2177 VGND.n26 VGND.n25 26.7302
R2178 VGND.n27 VGND.n26 26.7302
R2179 VGND.n1331 VGND.n27 26.7302
R2180 VGND.n31 VGND.n30 26.7302
R2181 VGND.n32 VGND.n31 26.7302
R2182 VGND.n1334 VGND.n32 26.7302
R2183 VGND.n1334 VGND.n35 26.7302
R2184 VGND.n37 VGND.n36 26.7302
R2185 VGND.n1337 VGND.n37 26.7302
R2186 VGND.n1337 VGND.n40 26.7302
R2187 VGND.n41 VGND.n40 26.7302
R2188 VGND.n1340 VGND.n42 26.7302
R2189 VGND.n1340 VGND.n45 26.7302
R2190 VGND.n46 VGND.n45 26.7302
R2191 VGND.n47 VGND.n46 26.7302
R2192 VGND.n1343 VGND.n50 26.7302
R2193 VGND.n51 VGND.n50 26.7302
R2194 VGND.n52 VGND.n51 26.7302
R2195 VGND.n1346 VGND.n52 26.7302
R2196 VGND.n56 VGND.n55 26.7302
R2197 VGND.n57 VGND.n56 26.7302
R2198 VGND.n1349 VGND.n57 26.7302
R2199 VGND.n1349 VGND.n60 26.7302
R2200 VGND.n62 VGND.n61 26.7302
R2201 VGND.n1352 VGND.n62 26.7302
R2202 VGND.n1352 VGND.n65 26.7302
R2203 VGND.n66 VGND.n65 26.7302
R2204 VGND.n1355 VGND.n67 26.7302
R2205 VGND.n1355 VGND.n70 26.7302
R2206 VGND.n71 VGND.n70 26.7302
R2207 VGND.n72 VGND.n71 26.7302
R2208 VGND.n1358 VGND.n75 26.7302
R2209 VGND.n76 VGND.n75 26.7302
R2210 VGND.n77 VGND.n76 26.7302
R2211 VGND.n1361 VGND.n77 26.7302
R2212 VGND.n81 VGND.n80 26.7302
R2213 VGND.n82 VGND.n81 26.7302
R2214 VGND.n1364 VGND.n82 26.7302
R2215 VGND.n1364 VGND.n85 26.7302
R2216 VGND.n87 VGND.n86 26.7302
R2217 VGND.n1367 VGND.n87 26.7302
R2218 VGND.n1367 VGND.n90 26.7302
R2219 VGND.n91 VGND.n90 26.7302
R2220 VGND.n632 VGND.n629 25.9877
R2221 VGND.n938 VGND.n630 25.9877
R2222 VGND.n937 VGND.n626 25.9877
R2223 VGND.n1300 VGND.t22 25.9877
R2224 VGND.n11 VGND.t27 25.9877
R2225 VGND.n103 VGND.n92 25.9877
R2226 VGND.n1561 VGND.n181 25.9877
R2227 VGND.n1566 VGND.n96 25.9877
R2228 VGND.n510 VGND.t1 25.2452
R2229 VGND.n17 VGND.t29 25.2452
R2230 VGND.n861 VGND.n625 24.9538
R2231 VGND.n1370 VGND.n101 24.9538
R2232 VGND.n1101 VGND.n627 24.9538
R2233 VGND.n1570 VGND.n93 24.9538
R2234 VGND.n1270 VGND.t26 24.5027
R2235 VGND.n1328 VGND.t16 24.5027
R2236 VGND.n530 VGND.t13 23.7602
R2237 VGND.t7 VGND.n30 23.7602
R2238 VGND.n1240 VGND.t30 23.0177
R2239 VGND.n36 VGND.t28 23.0177
R2240 VGND.n104 VGND.n102 22.7228
R2241 VGND.n1560 VGND.n407 22.7228
R2242 VGND.n408 VGND.n105 22.7228
R2243 VGND.n406 VGND.n404 22.7228
R2244 VGND.n405 VGND.n106 22.7228
R2245 VGND.n403 VGND.n401 22.7228
R2246 VGND.n402 VGND.n107 22.7228
R2247 VGND.n400 VGND.n398 22.7228
R2248 VGND.n399 VGND.n108 22.7228
R2249 VGND.n397 VGND.n395 22.7228
R2250 VGND.n396 VGND.n109 22.7228
R2251 VGND.n394 VGND.n392 22.7228
R2252 VGND.n393 VGND.n110 22.7228
R2253 VGND.n391 VGND.n389 22.7228
R2254 VGND.n390 VGND.n111 22.7228
R2255 VGND.n388 VGND.n386 22.7228
R2256 VGND.n387 VGND.n112 22.7228
R2257 VGND.n385 VGND.n383 22.7228
R2258 VGND.n384 VGND.n113 22.7228
R2259 VGND.n382 VGND.n380 22.7228
R2260 VGND.n381 VGND.n114 22.7228
R2261 VGND.n379 VGND.n377 22.7228
R2262 VGND.n378 VGND.n115 22.7228
R2263 VGND.n376 VGND.n374 22.7228
R2264 VGND.n375 VGND.n116 22.7228
R2265 VGND.n373 VGND.n371 22.7228
R2266 VGND.n372 VGND.n117 22.7228
R2267 VGND.n370 VGND.n368 22.7228
R2268 VGND.n369 VGND.n118 22.7228
R2269 VGND.n367 VGND.n365 22.7228
R2270 VGND.n366 VGND.n119 22.7228
R2271 VGND.n364 VGND.n362 22.7228
R2272 VGND.n363 VGND.n120 22.7228
R2273 VGND.n361 VGND.n359 22.7228
R2274 VGND.n360 VGND.n121 22.7228
R2275 VGND.n358 VGND.n356 22.7228
R2276 VGND.n357 VGND.n122 22.7228
R2277 VGND.n355 VGND.n353 22.7228
R2278 VGND.n354 VGND.n123 22.7228
R2279 VGND.n352 VGND.n350 22.7228
R2280 VGND.n351 VGND.n124 22.7228
R2281 VGND.n349 VGND.n347 22.7228
R2282 VGND.n348 VGND.n125 22.7228
R2283 VGND.n346 VGND.n344 22.7228
R2284 VGND.n345 VGND.n126 22.7228
R2285 VGND.n343 VGND.n341 22.7228
R2286 VGND.n342 VGND.n127 22.7228
R2287 VGND.n340 VGND.n338 22.7228
R2288 VGND.n339 VGND.n128 22.7228
R2289 VGND.n337 VGND.n335 22.7228
R2290 VGND.n336 VGND.n129 22.7228
R2291 VGND.n334 VGND.n332 22.7228
R2292 VGND.n333 VGND.n130 22.7228
R2293 VGND.n331 VGND.n329 22.7228
R2294 VGND.n330 VGND.n131 22.7228
R2295 VGND.n328 VGND.n326 22.7228
R2296 VGND.n327 VGND.n132 22.7228
R2297 VGND.n325 VGND.n323 22.7228
R2298 VGND.n324 VGND.n133 22.7228
R2299 VGND.n322 VGND.n320 22.7228
R2300 VGND.n321 VGND.n134 22.7228
R2301 VGND.n319 VGND.n317 22.7228
R2302 VGND.n318 VGND.n135 22.7228
R2303 VGND.n316 VGND.n314 22.7228
R2304 VGND.n315 VGND.n136 22.7228
R2305 VGND.n313 VGND.n311 22.7228
R2306 VGND.n312 VGND.n137 22.7228
R2307 VGND.n310 VGND.n308 22.7228
R2308 VGND.n309 VGND.n138 22.7228
R2309 VGND.n307 VGND.n305 22.7228
R2310 VGND.n306 VGND.n139 22.7228
R2311 VGND.n304 VGND.n302 22.7228
R2312 VGND.n303 VGND.n140 22.7228
R2313 VGND.n301 VGND.n299 22.7228
R2314 VGND.n300 VGND.n141 22.7228
R2315 VGND.n298 VGND.n296 22.7228
R2316 VGND.n297 VGND.n142 22.7228
R2317 VGND.n295 VGND.n293 22.7228
R2318 VGND.n294 VGND.n143 22.7228
R2319 VGND.n292 VGND.n290 22.7228
R2320 VGND.n291 VGND.n144 22.7228
R2321 VGND.n289 VGND.n287 22.7228
R2322 VGND.n288 VGND.n145 22.7228
R2323 VGND.n286 VGND.n284 22.7228
R2324 VGND.n285 VGND.n146 22.7228
R2325 VGND.n283 VGND.n281 22.7228
R2326 VGND.n282 VGND.n147 22.7228
R2327 VGND.n280 VGND.n278 22.7228
R2328 VGND.n279 VGND.n148 22.7228
R2329 VGND.n277 VGND.n275 22.7228
R2330 VGND.n276 VGND.n149 22.7228
R2331 VGND.n274 VGND.n272 22.7228
R2332 VGND.n273 VGND.n150 22.7228
R2333 VGND.n271 VGND.n269 22.7228
R2334 VGND.n270 VGND.n151 22.7228
R2335 VGND.n268 VGND.n266 22.7228
R2336 VGND.n267 VGND.n152 22.7228
R2337 VGND.n265 VGND.n263 22.7228
R2338 VGND.n264 VGND.n153 22.7228
R2339 VGND.n262 VGND.n260 22.7228
R2340 VGND.n261 VGND.n154 22.7228
R2341 VGND.n259 VGND.n257 22.7228
R2342 VGND.n258 VGND.n155 22.7228
R2343 VGND.n256 VGND.n254 22.7228
R2344 VGND.n255 VGND.n156 22.7228
R2345 VGND.n253 VGND.n251 22.7228
R2346 VGND.n252 VGND.n157 22.7228
R2347 VGND.n250 VGND.n248 22.7228
R2348 VGND.n249 VGND.n158 22.7228
R2349 VGND.n247 VGND.n245 22.7228
R2350 VGND.n246 VGND.n159 22.7228
R2351 VGND.n244 VGND.n242 22.7228
R2352 VGND.n243 VGND.n160 22.7228
R2353 VGND.n241 VGND.n239 22.7228
R2354 VGND.n240 VGND.n161 22.7228
R2355 VGND.n238 VGND.n236 22.7228
R2356 VGND.n237 VGND.n162 22.7228
R2357 VGND.n235 VGND.n233 22.7228
R2358 VGND.n234 VGND.n163 22.7228
R2359 VGND.n232 VGND.n230 22.7228
R2360 VGND.n231 VGND.n164 22.7228
R2361 VGND.n229 VGND.n227 22.7228
R2362 VGND.n228 VGND.n165 22.7228
R2363 VGND.n226 VGND.n224 22.7228
R2364 VGND.n225 VGND.n166 22.7228
R2365 VGND.n223 VGND.n221 22.7228
R2366 VGND.n222 VGND.n167 22.7228
R2367 VGND.n220 VGND.n218 22.7228
R2368 VGND.n219 VGND.n168 22.7228
R2369 VGND.n217 VGND.n215 22.7228
R2370 VGND.n216 VGND.n169 22.7228
R2371 VGND.n214 VGND.n212 22.7228
R2372 VGND.n213 VGND.n170 22.7228
R2373 VGND.n211 VGND.n209 22.7228
R2374 VGND.n210 VGND.n171 22.7228
R2375 VGND.n208 VGND.n206 22.7228
R2376 VGND.n207 VGND.n172 22.7228
R2377 VGND.n205 VGND.n203 22.7228
R2378 VGND.n204 VGND.n173 22.7228
R2379 VGND.n202 VGND.n200 22.7228
R2380 VGND.n201 VGND.n174 22.7228
R2381 VGND.n199 VGND.n197 22.7228
R2382 VGND.n198 VGND.n175 22.7228
R2383 VGND.n196 VGND.n194 22.7228
R2384 VGND.n195 VGND.n176 22.7228
R2385 VGND.n193 VGND.n191 22.7228
R2386 VGND.n192 VGND.n177 22.7228
R2387 VGND.n190 VGND.n188 22.7228
R2388 VGND.n189 VGND.n178 22.7228
R2389 VGND.n187 VGND.n185 22.7228
R2390 VGND.n186 VGND.n179 22.7228
R2391 VGND.n184 VGND.n182 22.7228
R2392 VGND.n183 VGND.n180 22.7228
R2393 VGND.n939 VGND.n633 22.7228
R2394 VGND.n859 VGND.n633 22.7228
R2395 VGND.n862 VGND.n634 22.7228
R2396 VGND.n857 VGND.n634 22.7228
R2397 VGND.n863 VGND.n635 22.7228
R2398 VGND.n855 VGND.n635 22.7228
R2399 VGND.n864 VGND.n636 22.7228
R2400 VGND.n853 VGND.n636 22.7228
R2401 VGND.n865 VGND.n637 22.7228
R2402 VGND.n851 VGND.n637 22.7228
R2403 VGND.n866 VGND.n638 22.7228
R2404 VGND.n849 VGND.n638 22.7228
R2405 VGND.n867 VGND.n639 22.7228
R2406 VGND.n847 VGND.n639 22.7228
R2407 VGND.n868 VGND.n640 22.7228
R2408 VGND.n845 VGND.n640 22.7228
R2409 VGND.n869 VGND.n641 22.7228
R2410 VGND.n843 VGND.n641 22.7228
R2411 VGND.n870 VGND.n642 22.7228
R2412 VGND.n841 VGND.n642 22.7228
R2413 VGND.n871 VGND.n643 22.7228
R2414 VGND.n839 VGND.n643 22.7228
R2415 VGND.n872 VGND.n644 22.7228
R2416 VGND.n837 VGND.n644 22.7228
R2417 VGND.n873 VGND.n645 22.7228
R2418 VGND.n835 VGND.n645 22.7228
R2419 VGND.n874 VGND.n646 22.7228
R2420 VGND.n833 VGND.n646 22.7228
R2421 VGND.n875 VGND.n647 22.7228
R2422 VGND.n831 VGND.n647 22.7228
R2423 VGND.n876 VGND.n648 22.7228
R2424 VGND.n829 VGND.n648 22.7228
R2425 VGND.n877 VGND.n649 22.7228
R2426 VGND.n827 VGND.n649 22.7228
R2427 VGND.n878 VGND.n650 22.7228
R2428 VGND.n825 VGND.n650 22.7228
R2429 VGND.n879 VGND.n651 22.7228
R2430 VGND.n823 VGND.n651 22.7228
R2431 VGND.n880 VGND.n652 22.7228
R2432 VGND.n821 VGND.n652 22.7228
R2433 VGND.n881 VGND.n653 22.7228
R2434 VGND.n819 VGND.n653 22.7228
R2435 VGND.n882 VGND.n654 22.7228
R2436 VGND.n817 VGND.n654 22.7228
R2437 VGND.n883 VGND.n655 22.7228
R2438 VGND.n815 VGND.n655 22.7228
R2439 VGND.n884 VGND.n656 22.7228
R2440 VGND.n813 VGND.n656 22.7228
R2441 VGND.n885 VGND.n657 22.7228
R2442 VGND.n811 VGND.n657 22.7228
R2443 VGND.n886 VGND.n658 22.7228
R2444 VGND.n809 VGND.n658 22.7228
R2445 VGND.n887 VGND.n659 22.7228
R2446 VGND.n807 VGND.n659 22.7228
R2447 VGND.n888 VGND.n660 22.7228
R2448 VGND.n805 VGND.n660 22.7228
R2449 VGND.n889 VGND.n661 22.7228
R2450 VGND.n803 VGND.n661 22.7228
R2451 VGND.n890 VGND.n662 22.7228
R2452 VGND.n801 VGND.n662 22.7228
R2453 VGND.n891 VGND.n663 22.7228
R2454 VGND.n799 VGND.n663 22.7228
R2455 VGND.n892 VGND.n664 22.7228
R2456 VGND.n797 VGND.n664 22.7228
R2457 VGND.n893 VGND.n665 22.7228
R2458 VGND.n795 VGND.n665 22.7228
R2459 VGND.n894 VGND.n666 22.7228
R2460 VGND.n793 VGND.n666 22.7228
R2461 VGND.n895 VGND.n667 22.7228
R2462 VGND.n791 VGND.n667 22.7228
R2463 VGND.n896 VGND.n668 22.7228
R2464 VGND.n789 VGND.n668 22.7228
R2465 VGND.n897 VGND.n669 22.7228
R2466 VGND.n787 VGND.n669 22.7228
R2467 VGND.n898 VGND.n670 22.7228
R2468 VGND.n785 VGND.n670 22.7228
R2469 VGND.n899 VGND.n671 22.7228
R2470 VGND.n783 VGND.n671 22.7228
R2471 VGND.n900 VGND.n672 22.7228
R2472 VGND.n781 VGND.n672 22.7228
R2473 VGND.n901 VGND.n673 22.7228
R2474 VGND.n779 VGND.n673 22.7228
R2475 VGND.n902 VGND.n674 22.7228
R2476 VGND.n777 VGND.n674 22.7228
R2477 VGND.n903 VGND.n675 22.7228
R2478 VGND.n775 VGND.n675 22.7228
R2479 VGND.n904 VGND.n676 22.7228
R2480 VGND.n773 VGND.n676 22.7228
R2481 VGND.n905 VGND.n677 22.7228
R2482 VGND.n771 VGND.n677 22.7228
R2483 VGND.n906 VGND.n678 22.7228
R2484 VGND.n769 VGND.n678 22.7228
R2485 VGND.n907 VGND.n679 22.7228
R2486 VGND.n767 VGND.n679 22.7228
R2487 VGND.n908 VGND.n680 22.7228
R2488 VGND.n765 VGND.n680 22.7228
R2489 VGND.n909 VGND.n681 22.7228
R2490 VGND.n763 VGND.n681 22.7228
R2491 VGND.n910 VGND.n682 22.7228
R2492 VGND.n761 VGND.n682 22.7228
R2493 VGND.n911 VGND.n683 22.7228
R2494 VGND.n759 VGND.n683 22.7228
R2495 VGND.n912 VGND.n684 22.7228
R2496 VGND.n757 VGND.n684 22.7228
R2497 VGND.n913 VGND.n685 22.7228
R2498 VGND.n755 VGND.n685 22.7228
R2499 VGND.n914 VGND.n686 22.7228
R2500 VGND.n753 VGND.n686 22.7228
R2501 VGND.n915 VGND.n687 22.7228
R2502 VGND.n751 VGND.n687 22.7228
R2503 VGND.n916 VGND.n688 22.7228
R2504 VGND.n749 VGND.n688 22.7228
R2505 VGND.n917 VGND.n689 22.7228
R2506 VGND.n747 VGND.n689 22.7228
R2507 VGND.n918 VGND.n690 22.7228
R2508 VGND.n745 VGND.n690 22.7228
R2509 VGND.n919 VGND.n691 22.7228
R2510 VGND.n743 VGND.n691 22.7228
R2511 VGND.n920 VGND.n692 22.7228
R2512 VGND.n741 VGND.n692 22.7228
R2513 VGND.n921 VGND.n693 22.7228
R2514 VGND.n739 VGND.n693 22.7228
R2515 VGND.n922 VGND.n694 22.7228
R2516 VGND.n737 VGND.n694 22.7228
R2517 VGND.n923 VGND.n695 22.7228
R2518 VGND.n735 VGND.n695 22.7228
R2519 VGND.n924 VGND.n696 22.7228
R2520 VGND.n733 VGND.n696 22.7228
R2521 VGND.n925 VGND.n697 22.7228
R2522 VGND.n731 VGND.n697 22.7228
R2523 VGND.n926 VGND.n698 22.7228
R2524 VGND.n729 VGND.n698 22.7228
R2525 VGND.n927 VGND.n699 22.7228
R2526 VGND.n727 VGND.n699 22.7228
R2527 VGND.n928 VGND.n700 22.7228
R2528 VGND.n725 VGND.n700 22.7228
R2529 VGND.n929 VGND.n701 22.7228
R2530 VGND.n723 VGND.n701 22.7228
R2531 VGND.n930 VGND.n702 22.7228
R2532 VGND.n721 VGND.n702 22.7228
R2533 VGND.n931 VGND.n703 22.7228
R2534 VGND.n719 VGND.n703 22.7228
R2535 VGND.n932 VGND.n704 22.7228
R2536 VGND.n717 VGND.n704 22.7228
R2537 VGND.n933 VGND.n705 22.7228
R2538 VGND.n715 VGND.n705 22.7228
R2539 VGND.n934 VGND.n706 22.7228
R2540 VGND.n713 VGND.n706 22.7228
R2541 VGND.n935 VGND.n707 22.7228
R2542 VGND.n711 VGND.n707 22.7228
R2543 VGND.n936 VGND.n708 22.7228
R2544 VGND.n709 VGND.n708 22.7228
R2545 VGND.n1100 VGND.n631 22.7228
R2546 VGND.n1098 VGND.n939 22.7228
R2547 VGND.n860 VGND.n859 22.7228
R2548 VGND.n862 VGND.n860 22.7228
R2549 VGND.n858 VGND.n857 22.7228
R2550 VGND.n863 VGND.n858 22.7228
R2551 VGND.n856 VGND.n855 22.7228
R2552 VGND.n864 VGND.n856 22.7228
R2553 VGND.n854 VGND.n853 22.7228
R2554 VGND.n865 VGND.n854 22.7228
R2555 VGND.n852 VGND.n851 22.7228
R2556 VGND.n866 VGND.n852 22.7228
R2557 VGND.n850 VGND.n849 22.7228
R2558 VGND.n867 VGND.n850 22.7228
R2559 VGND.n848 VGND.n847 22.7228
R2560 VGND.n868 VGND.n848 22.7228
R2561 VGND.n846 VGND.n845 22.7228
R2562 VGND.n869 VGND.n846 22.7228
R2563 VGND.n844 VGND.n843 22.7228
R2564 VGND.n870 VGND.n844 22.7228
R2565 VGND.n842 VGND.n841 22.7228
R2566 VGND.n871 VGND.n842 22.7228
R2567 VGND.n840 VGND.n839 22.7228
R2568 VGND.n872 VGND.n840 22.7228
R2569 VGND.n838 VGND.n837 22.7228
R2570 VGND.n873 VGND.n838 22.7228
R2571 VGND.n836 VGND.n835 22.7228
R2572 VGND.n874 VGND.n836 22.7228
R2573 VGND.n834 VGND.n833 22.7228
R2574 VGND.n875 VGND.n834 22.7228
R2575 VGND.n832 VGND.n831 22.7228
R2576 VGND.n876 VGND.n832 22.7228
R2577 VGND.n830 VGND.n829 22.7228
R2578 VGND.n877 VGND.n830 22.7228
R2579 VGND.n828 VGND.n827 22.7228
R2580 VGND.n878 VGND.n828 22.7228
R2581 VGND.n826 VGND.n825 22.7228
R2582 VGND.n879 VGND.n826 22.7228
R2583 VGND.n824 VGND.n823 22.7228
R2584 VGND.n880 VGND.n824 22.7228
R2585 VGND.n822 VGND.n821 22.7228
R2586 VGND.n881 VGND.n822 22.7228
R2587 VGND.n820 VGND.n819 22.7228
R2588 VGND.n882 VGND.n820 22.7228
R2589 VGND.n818 VGND.n817 22.7228
R2590 VGND.n883 VGND.n818 22.7228
R2591 VGND.n816 VGND.n815 22.7228
R2592 VGND.n884 VGND.n816 22.7228
R2593 VGND.n814 VGND.n813 22.7228
R2594 VGND.n885 VGND.n814 22.7228
R2595 VGND.n812 VGND.n811 22.7228
R2596 VGND.n886 VGND.n812 22.7228
R2597 VGND.n810 VGND.n809 22.7228
R2598 VGND.n887 VGND.n810 22.7228
R2599 VGND.n808 VGND.n807 22.7228
R2600 VGND.n888 VGND.n808 22.7228
R2601 VGND.n806 VGND.n805 22.7228
R2602 VGND.n889 VGND.n806 22.7228
R2603 VGND.n804 VGND.n803 22.7228
R2604 VGND.n890 VGND.n804 22.7228
R2605 VGND.n802 VGND.n801 22.7228
R2606 VGND.n891 VGND.n802 22.7228
R2607 VGND.n800 VGND.n799 22.7228
R2608 VGND.n892 VGND.n800 22.7228
R2609 VGND.n798 VGND.n797 22.7228
R2610 VGND.n893 VGND.n798 22.7228
R2611 VGND.n796 VGND.n795 22.7228
R2612 VGND.n894 VGND.n796 22.7228
R2613 VGND.n794 VGND.n793 22.7228
R2614 VGND.n895 VGND.n794 22.7228
R2615 VGND.n792 VGND.n791 22.7228
R2616 VGND.n896 VGND.n792 22.7228
R2617 VGND.n790 VGND.n789 22.7228
R2618 VGND.n897 VGND.n790 22.7228
R2619 VGND.n788 VGND.n787 22.7228
R2620 VGND.n898 VGND.n788 22.7228
R2621 VGND.n786 VGND.n785 22.7228
R2622 VGND.n899 VGND.n786 22.7228
R2623 VGND.n784 VGND.n783 22.7228
R2624 VGND.n900 VGND.n784 22.7228
R2625 VGND.n782 VGND.n781 22.7228
R2626 VGND.n901 VGND.n782 22.7228
R2627 VGND.n780 VGND.n779 22.7228
R2628 VGND.n902 VGND.n780 22.7228
R2629 VGND.n778 VGND.n777 22.7228
R2630 VGND.n903 VGND.n778 22.7228
R2631 VGND.n776 VGND.n775 22.7228
R2632 VGND.n904 VGND.n776 22.7228
R2633 VGND.n774 VGND.n773 22.7228
R2634 VGND.n905 VGND.n774 22.7228
R2635 VGND.n772 VGND.n771 22.7228
R2636 VGND.n906 VGND.n772 22.7228
R2637 VGND.n770 VGND.n769 22.7228
R2638 VGND.n907 VGND.n770 22.7228
R2639 VGND.n768 VGND.n767 22.7228
R2640 VGND.n908 VGND.n768 22.7228
R2641 VGND.n766 VGND.n765 22.7228
R2642 VGND.n909 VGND.n766 22.7228
R2643 VGND.n764 VGND.n763 22.7228
R2644 VGND.n910 VGND.n764 22.7228
R2645 VGND.n762 VGND.n761 22.7228
R2646 VGND.n911 VGND.n762 22.7228
R2647 VGND.n760 VGND.n759 22.7228
R2648 VGND.n912 VGND.n760 22.7228
R2649 VGND.n758 VGND.n757 22.7228
R2650 VGND.n913 VGND.n758 22.7228
R2651 VGND.n756 VGND.n755 22.7228
R2652 VGND.n914 VGND.n756 22.7228
R2653 VGND.n754 VGND.n753 22.7228
R2654 VGND.n915 VGND.n754 22.7228
R2655 VGND.n752 VGND.n751 22.7228
R2656 VGND.n916 VGND.n752 22.7228
R2657 VGND.n750 VGND.n749 22.7228
R2658 VGND.n917 VGND.n750 22.7228
R2659 VGND.n748 VGND.n747 22.7228
R2660 VGND.n918 VGND.n748 22.7228
R2661 VGND.n746 VGND.n745 22.7228
R2662 VGND.n919 VGND.n746 22.7228
R2663 VGND.n744 VGND.n743 22.7228
R2664 VGND.n920 VGND.n744 22.7228
R2665 VGND.n742 VGND.n741 22.7228
R2666 VGND.n921 VGND.n742 22.7228
R2667 VGND.n740 VGND.n739 22.7228
R2668 VGND.n922 VGND.n740 22.7228
R2669 VGND.n738 VGND.n737 22.7228
R2670 VGND.n923 VGND.n738 22.7228
R2671 VGND.n736 VGND.n735 22.7228
R2672 VGND.n924 VGND.n736 22.7228
R2673 VGND.n734 VGND.n733 22.7228
R2674 VGND.n925 VGND.n734 22.7228
R2675 VGND.n732 VGND.n731 22.7228
R2676 VGND.n926 VGND.n732 22.7228
R2677 VGND.n730 VGND.n729 22.7228
R2678 VGND.n927 VGND.n730 22.7228
R2679 VGND.n728 VGND.n727 22.7228
R2680 VGND.n928 VGND.n728 22.7228
R2681 VGND.n726 VGND.n725 22.7228
R2682 VGND.n929 VGND.n726 22.7228
R2683 VGND.n724 VGND.n723 22.7228
R2684 VGND.n930 VGND.n724 22.7228
R2685 VGND.n722 VGND.n721 22.7228
R2686 VGND.n931 VGND.n722 22.7228
R2687 VGND.n720 VGND.n719 22.7228
R2688 VGND.n932 VGND.n720 22.7228
R2689 VGND.n718 VGND.n717 22.7228
R2690 VGND.n933 VGND.n718 22.7228
R2691 VGND.n716 VGND.n715 22.7228
R2692 VGND.n934 VGND.n716 22.7228
R2693 VGND.n714 VGND.n713 22.7228
R2694 VGND.n935 VGND.n714 22.7228
R2695 VGND.n712 VGND.n711 22.7228
R2696 VGND.n936 VGND.n712 22.7228
R2697 VGND.n710 VGND.n709 22.7228
R2698 VGND.n710 VGND.n631 22.7228
R2699 VGND.n184 VGND.n183 22.7228
R2700 VGND.n182 VGND.n179 22.7228
R2701 VGND.n187 VGND.n186 22.7228
R2702 VGND.n185 VGND.n178 22.7228
R2703 VGND.n190 VGND.n189 22.7228
R2704 VGND.n188 VGND.n177 22.7228
R2705 VGND.n193 VGND.n192 22.7228
R2706 VGND.n191 VGND.n176 22.7228
R2707 VGND.n196 VGND.n195 22.7228
R2708 VGND.n194 VGND.n175 22.7228
R2709 VGND.n199 VGND.n198 22.7228
R2710 VGND.n197 VGND.n174 22.7228
R2711 VGND.n202 VGND.n201 22.7228
R2712 VGND.n200 VGND.n173 22.7228
R2713 VGND.n205 VGND.n204 22.7228
R2714 VGND.n203 VGND.n172 22.7228
R2715 VGND.n208 VGND.n207 22.7228
R2716 VGND.n206 VGND.n171 22.7228
R2717 VGND.n211 VGND.n210 22.7228
R2718 VGND.n209 VGND.n170 22.7228
R2719 VGND.n214 VGND.n213 22.7228
R2720 VGND.n212 VGND.n169 22.7228
R2721 VGND.n217 VGND.n216 22.7228
R2722 VGND.n215 VGND.n168 22.7228
R2723 VGND.n220 VGND.n219 22.7228
R2724 VGND.n218 VGND.n167 22.7228
R2725 VGND.n223 VGND.n222 22.7228
R2726 VGND.n221 VGND.n166 22.7228
R2727 VGND.n226 VGND.n225 22.7228
R2728 VGND.n224 VGND.n165 22.7228
R2729 VGND.n229 VGND.n228 22.7228
R2730 VGND.n227 VGND.n164 22.7228
R2731 VGND.n232 VGND.n231 22.7228
R2732 VGND.n230 VGND.n163 22.7228
R2733 VGND.n235 VGND.n234 22.7228
R2734 VGND.n233 VGND.n162 22.7228
R2735 VGND.n238 VGND.n237 22.7228
R2736 VGND.n236 VGND.n161 22.7228
R2737 VGND.n241 VGND.n240 22.7228
R2738 VGND.n239 VGND.n160 22.7228
R2739 VGND.n244 VGND.n243 22.7228
R2740 VGND.n242 VGND.n159 22.7228
R2741 VGND.n247 VGND.n246 22.7228
R2742 VGND.n245 VGND.n158 22.7228
R2743 VGND.n250 VGND.n249 22.7228
R2744 VGND.n248 VGND.n157 22.7228
R2745 VGND.n253 VGND.n252 22.7228
R2746 VGND.n251 VGND.n156 22.7228
R2747 VGND.n256 VGND.n255 22.7228
R2748 VGND.n254 VGND.n155 22.7228
R2749 VGND.n259 VGND.n258 22.7228
R2750 VGND.n257 VGND.n154 22.7228
R2751 VGND.n262 VGND.n261 22.7228
R2752 VGND.n260 VGND.n153 22.7228
R2753 VGND.n265 VGND.n264 22.7228
R2754 VGND.n263 VGND.n152 22.7228
R2755 VGND.n268 VGND.n267 22.7228
R2756 VGND.n266 VGND.n151 22.7228
R2757 VGND.n271 VGND.n270 22.7228
R2758 VGND.n269 VGND.n150 22.7228
R2759 VGND.n274 VGND.n273 22.7228
R2760 VGND.n272 VGND.n149 22.7228
R2761 VGND.n277 VGND.n276 22.7228
R2762 VGND.n275 VGND.n148 22.7228
R2763 VGND.n280 VGND.n279 22.7228
R2764 VGND.n278 VGND.n147 22.7228
R2765 VGND.n283 VGND.n282 22.7228
R2766 VGND.n281 VGND.n146 22.7228
R2767 VGND.n286 VGND.n285 22.7228
R2768 VGND.n284 VGND.n145 22.7228
R2769 VGND.n289 VGND.n288 22.7228
R2770 VGND.n287 VGND.n144 22.7228
R2771 VGND.n292 VGND.n291 22.7228
R2772 VGND.n290 VGND.n143 22.7228
R2773 VGND.n295 VGND.n294 22.7228
R2774 VGND.n293 VGND.n142 22.7228
R2775 VGND.n298 VGND.n297 22.7228
R2776 VGND.n296 VGND.n141 22.7228
R2777 VGND.n301 VGND.n300 22.7228
R2778 VGND.n299 VGND.n140 22.7228
R2779 VGND.n304 VGND.n303 22.7228
R2780 VGND.n302 VGND.n139 22.7228
R2781 VGND.n307 VGND.n306 22.7228
R2782 VGND.n305 VGND.n138 22.7228
R2783 VGND.n310 VGND.n309 22.7228
R2784 VGND.n308 VGND.n137 22.7228
R2785 VGND.n313 VGND.n312 22.7228
R2786 VGND.n311 VGND.n136 22.7228
R2787 VGND.n316 VGND.n315 22.7228
R2788 VGND.n314 VGND.n135 22.7228
R2789 VGND.n319 VGND.n318 22.7228
R2790 VGND.n317 VGND.n134 22.7228
R2791 VGND.n322 VGND.n321 22.7228
R2792 VGND.n320 VGND.n133 22.7228
R2793 VGND.n325 VGND.n324 22.7228
R2794 VGND.n323 VGND.n132 22.7228
R2795 VGND.n328 VGND.n327 22.7228
R2796 VGND.n326 VGND.n131 22.7228
R2797 VGND.n331 VGND.n330 22.7228
R2798 VGND.n329 VGND.n130 22.7228
R2799 VGND.n334 VGND.n333 22.7228
R2800 VGND.n332 VGND.n129 22.7228
R2801 VGND.n337 VGND.n336 22.7228
R2802 VGND.n335 VGND.n128 22.7228
R2803 VGND.n340 VGND.n339 22.7228
R2804 VGND.n338 VGND.n127 22.7228
R2805 VGND.n343 VGND.n342 22.7228
R2806 VGND.n341 VGND.n126 22.7228
R2807 VGND.n346 VGND.n345 22.7228
R2808 VGND.n344 VGND.n125 22.7228
R2809 VGND.n349 VGND.n348 22.7228
R2810 VGND.n347 VGND.n124 22.7228
R2811 VGND.n352 VGND.n351 22.7228
R2812 VGND.n350 VGND.n123 22.7228
R2813 VGND.n355 VGND.n354 22.7228
R2814 VGND.n353 VGND.n122 22.7228
R2815 VGND.n358 VGND.n357 22.7228
R2816 VGND.n356 VGND.n121 22.7228
R2817 VGND.n361 VGND.n360 22.7228
R2818 VGND.n359 VGND.n120 22.7228
R2819 VGND.n364 VGND.n363 22.7228
R2820 VGND.n362 VGND.n119 22.7228
R2821 VGND.n367 VGND.n366 22.7228
R2822 VGND.n365 VGND.n118 22.7228
R2823 VGND.n370 VGND.n369 22.7228
R2824 VGND.n368 VGND.n117 22.7228
R2825 VGND.n373 VGND.n372 22.7228
R2826 VGND.n371 VGND.n116 22.7228
R2827 VGND.n376 VGND.n375 22.7228
R2828 VGND.n374 VGND.n115 22.7228
R2829 VGND.n379 VGND.n378 22.7228
R2830 VGND.n377 VGND.n114 22.7228
R2831 VGND.n382 VGND.n381 22.7228
R2832 VGND.n380 VGND.n113 22.7228
R2833 VGND.n385 VGND.n384 22.7228
R2834 VGND.n383 VGND.n112 22.7228
R2835 VGND.n388 VGND.n387 22.7228
R2836 VGND.n386 VGND.n111 22.7228
R2837 VGND.n391 VGND.n390 22.7228
R2838 VGND.n389 VGND.n110 22.7228
R2839 VGND.n394 VGND.n393 22.7228
R2840 VGND.n392 VGND.n109 22.7228
R2841 VGND.n397 VGND.n396 22.7228
R2842 VGND.n395 VGND.n108 22.7228
R2843 VGND.n400 VGND.n399 22.7228
R2844 VGND.n398 VGND.n107 22.7228
R2845 VGND.n403 VGND.n402 22.7228
R2846 VGND.n401 VGND.n106 22.7228
R2847 VGND.n406 VGND.n405 22.7228
R2848 VGND.n404 VGND.n105 22.7228
R2849 VGND.n1560 VGND.n408 22.7228
R2850 VGND.n407 VGND.n104 22.7228
R2851 VGND.n1562 VGND.n102 22.7228
R2852 VGND.n940 VGND.n861 22.3272
R2853 VGND.n101 VGND.n98 22.3272
R2854 VGND.n1102 VGND.n1101 22.3272
R2855 VGND.n95 VGND.n93 22.3272
R2856 VGND.n550 VGND.t3 22.2752
R2857 VGND.n42 VGND.t19 22.2752
R2858 VGND.n1210 VGND.t4 21.5327
R2859 VGND.n1343 VGND.t11 21.5327
R2860 VGND.n570 VGND.t2 20.7902
R2861 VGND.t20 VGND.n55 20.7902
R2862 VGND.n941 VGND.n940 20.1701
R2863 VGND.n1567 VGND.n95 20.1701
R2864 VGND.n1565 VGND.n98 20.1692
R2865 VGND.n1103 VGND.n1102 20.1692
R2866 VGND.n1180 VGND.t14 20.0478
R2867 VGND.n61 VGND.t17 20.0478
R2868 VGND.n590 VGND.t0 19.3053
R2869 VGND.n67 VGND.t12 19.3053
R2870 VGND.n1150 VGND.t6 18.5628
R2871 VGND.n1358 VGND.t31 18.5628
R2872 VGND.n610 VGND.t21 17.8203
R2873 VGND.t5 VGND.n80 17.8203
R2874 VGND.n1120 VGND.t8 17.0778
R2875 VGND.n86 VGND.t23 17.0778
R2876 VGND.t8 VGND.n614 9.65288
R2877 VGND.t23 VGND.n85 9.65288
R2878 VGND.n1138 VGND.t21 8.91039
R2879 VGND.n1361 VGND.t5 8.91039
R2880 VGND.t6 VGND.n594 8.1679
R2881 VGND.t31 VGND.n72 8.1679
R2882 VGND.n1168 VGND.t0 7.42541
R2883 VGND.t12 VGND.n66 7.42541
R2884 VGND.t14 VGND.n574 6.68292
R2885 VGND.t17 VGND.n60 6.68292
R2886 VGND.n1198 VGND.t2 5.94043
R2887 VGND.n1346 VGND.t20 5.94043
R2888 VGND.t4 VGND.n554 5.19793
R2889 VGND.t11 VGND.n47 5.19793
R2890 VGND.n1479 VGND 4.59467
R2891 VGND.n1228 VGND.t3 4.45544
R2892 VGND.t19 VGND.n41 4.45544
R2893 VGND.n1097 VGND.n942 3.92583
R2894 VGND.n1104 VGND.n628 3.92583
R2895 VGND.n1564 VGND.n1563 3.92583
R2896 VGND.n1568 VGND.n94 3.92583
R2897 VGND.t30 VGND.n534 3.71295
R2898 VGND.t28 VGND.n35 3.71295
R2899 VGND.n1097 VGND.n1096 3.0725
R2900 VGND.n1096 VGND.n1095 3.0725
R2901 VGND.n1095 VGND.n1094 3.0725
R2902 VGND.n1094 VGND.n1093 3.0725
R2903 VGND.n1093 VGND.n1092 3.0725
R2904 VGND.n1092 VGND.n1091 3.0725
R2905 VGND.n1091 VGND.n1090 3.0725
R2906 VGND.n1090 VGND.n1089 3.0725
R2907 VGND.n1089 VGND.n1088 3.0725
R2908 VGND.n1088 VGND.n1087 3.0725
R2909 VGND.n1087 VGND.n1086 3.0725
R2910 VGND.n1086 VGND.n1085 3.0725
R2911 VGND.n1085 VGND.n1084 3.0725
R2912 VGND.n1084 VGND.n1083 3.0725
R2913 VGND.n1083 VGND.n1082 3.0725
R2914 VGND.n1082 VGND.n1081 3.0725
R2915 VGND.n1081 VGND.n1080 3.0725
R2916 VGND.n1080 VGND.n1079 3.0725
R2917 VGND.n1079 VGND.n1078 3.0725
R2918 VGND.n1078 VGND.n1077 3.0725
R2919 VGND.n1077 VGND.n1076 3.0725
R2920 VGND.n1076 VGND.n1075 3.0725
R2921 VGND.n1075 VGND.n1074 3.0725
R2922 VGND.n1074 VGND.n1073 3.0725
R2923 VGND.n1073 VGND.n1072 3.0725
R2924 VGND.n1072 VGND.n1071 3.0725
R2925 VGND.n1071 VGND.n1070 3.0725
R2926 VGND.n1070 VGND.n1069 3.0725
R2927 VGND.n1069 VGND.n1068 3.0725
R2928 VGND.n1068 VGND.n1067 3.0725
R2929 VGND.n1067 VGND.n1066 3.0725
R2930 VGND.n1066 VGND.n1065 3.0725
R2931 VGND.n1065 VGND.n1064 3.0725
R2932 VGND.n1064 VGND.n1063 3.0725
R2933 VGND.n1063 VGND.n1062 3.0725
R2934 VGND.n1062 VGND.n1061 3.0725
R2935 VGND.n1061 VGND.n1060 3.0725
R2936 VGND.n1060 VGND.n1059 3.0725
R2937 VGND.n1059 VGND.n1058 3.0725
R2938 VGND.n1058 VGND.n1057 3.0725
R2939 VGND.n1057 VGND.n1056 3.0725
R2940 VGND.n1056 VGND.n1055 3.0725
R2941 VGND.n1055 VGND.n1054 3.0725
R2942 VGND.n1054 VGND.n1053 3.0725
R2943 VGND.n1053 VGND.n1052 3.0725
R2944 VGND.n1052 VGND.n1051 3.0725
R2945 VGND.n1051 VGND.n1050 3.0725
R2946 VGND.n1050 VGND.n1049 3.0725
R2947 VGND.n1049 VGND.n1048 3.0725
R2948 VGND.n1048 VGND.n1047 3.0725
R2949 VGND.n1047 VGND.n1046 3.0725
R2950 VGND.n1046 VGND.n1045 3.0725
R2951 VGND.n1045 VGND.n1044 3.0725
R2952 VGND.n1044 VGND.n1043 3.0725
R2953 VGND.n1043 VGND.n1042 3.0725
R2954 VGND.n1042 VGND.n1041 3.0725
R2955 VGND.n1041 VGND.n1040 3.0725
R2956 VGND.n1040 VGND.n1039 3.0725
R2957 VGND.n1039 VGND.n1038 3.0725
R2958 VGND.n1038 VGND.n1037 3.0725
R2959 VGND.n1037 VGND.n1036 3.0725
R2960 VGND.n1036 VGND.n1035 3.0725
R2961 VGND.n1035 VGND.n1034 3.0725
R2962 VGND.n1034 VGND.n1033 3.0725
R2963 VGND.n1033 VGND.n1032 3.0725
R2964 VGND.n1032 VGND.n1031 3.0725
R2965 VGND.n1031 VGND.n1030 3.0725
R2966 VGND.n1030 VGND.n1029 3.0725
R2967 VGND.n1029 VGND.n1028 3.0725
R2968 VGND.n1028 VGND.n1027 3.0725
R2969 VGND.n1027 VGND.n1026 3.0725
R2970 VGND.n1026 VGND.n1025 3.0725
R2971 VGND.n1025 VGND.n1024 3.0725
R2972 VGND.n1024 VGND.n1023 3.0725
R2973 VGND.n1023 VGND.n1022 3.0725
R2974 VGND.n1022 VGND.n1021 3.0725
R2975 VGND.n1018 VGND.n1017 3.0725
R2976 VGND.n1017 VGND.n1016 3.0725
R2977 VGND.n1016 VGND.n1015 3.0725
R2978 VGND.n1015 VGND.n1014 3.0725
R2979 VGND.n1014 VGND.n1013 3.0725
R2980 VGND.n1013 VGND.n1012 3.0725
R2981 VGND.n1012 VGND.n1011 3.0725
R2982 VGND.n1011 VGND.n1010 3.0725
R2983 VGND.n1010 VGND.n1009 3.0725
R2984 VGND.n1009 VGND.n1008 3.0725
R2985 VGND.n1008 VGND.n1007 3.0725
R2986 VGND.n1007 VGND.n1006 3.0725
R2987 VGND.n1006 VGND.n1005 3.0725
R2988 VGND.n1005 VGND.n1004 3.0725
R2989 VGND.n1004 VGND.n1003 3.0725
R2990 VGND.n1003 VGND.n1002 3.0725
R2991 VGND.n1002 VGND.n1001 3.0725
R2992 VGND.n1001 VGND.n1000 3.0725
R2993 VGND.n1000 VGND.n999 3.0725
R2994 VGND.n999 VGND.n998 3.0725
R2995 VGND.n998 VGND.n997 3.0725
R2996 VGND.n997 VGND.n996 3.0725
R2997 VGND.n996 VGND.n995 3.0725
R2998 VGND.n995 VGND.n994 3.0725
R2999 VGND.n994 VGND.n993 3.0725
R3000 VGND.n993 VGND.n992 3.0725
R3001 VGND.n992 VGND.n991 3.0725
R3002 VGND.n991 VGND.n990 3.0725
R3003 VGND.n990 VGND.n989 3.0725
R3004 VGND.n989 VGND.n988 3.0725
R3005 VGND.n988 VGND.n987 3.0725
R3006 VGND.n987 VGND.n986 3.0725
R3007 VGND.n986 VGND.n985 3.0725
R3008 VGND.n985 VGND.n984 3.0725
R3009 VGND.n984 VGND.n983 3.0725
R3010 VGND.n983 VGND.n982 3.0725
R3011 VGND.n982 VGND.n981 3.0725
R3012 VGND.n981 VGND.n980 3.0725
R3013 VGND.n980 VGND.n979 3.0725
R3014 VGND.n979 VGND.n978 3.0725
R3015 VGND.n978 VGND.n977 3.0725
R3016 VGND.n977 VGND.n976 3.0725
R3017 VGND.n976 VGND.n975 3.0725
R3018 VGND.n975 VGND.n974 3.0725
R3019 VGND.n974 VGND.n973 3.0725
R3020 VGND.n973 VGND.n972 3.0725
R3021 VGND.n972 VGND.n971 3.0725
R3022 VGND.n971 VGND.n970 3.0725
R3023 VGND.n970 VGND.n969 3.0725
R3024 VGND.n969 VGND.n968 3.0725
R3025 VGND.n968 VGND.n967 3.0725
R3026 VGND.n967 VGND.n966 3.0725
R3027 VGND.n966 VGND.n965 3.0725
R3028 VGND.n965 VGND.n964 3.0725
R3029 VGND.n964 VGND.n963 3.0725
R3030 VGND.n963 VGND.n962 3.0725
R3031 VGND.n962 VGND.n961 3.0725
R3032 VGND.n961 VGND.n960 3.0725
R3033 VGND.n960 VGND.n959 3.0725
R3034 VGND.n959 VGND.n958 3.0725
R3035 VGND.n958 VGND.n957 3.0725
R3036 VGND.n957 VGND.n956 3.0725
R3037 VGND.n956 VGND.n955 3.0725
R3038 VGND.n955 VGND.n954 3.0725
R3039 VGND.n954 VGND.n953 3.0725
R3040 VGND.n953 VGND.n952 3.0725
R3041 VGND.n952 VGND.n951 3.0725
R3042 VGND.n951 VGND.n950 3.0725
R3043 VGND.n950 VGND.n949 3.0725
R3044 VGND.n949 VGND.n948 3.0725
R3045 VGND.n948 VGND.n947 3.0725
R3046 VGND.n947 VGND.n946 3.0725
R3047 VGND.n946 VGND.n945 3.0725
R3048 VGND.n945 VGND.n944 3.0725
R3049 VGND.n944 VGND.n943 3.0725
R3050 VGND.n943 VGND.n628 3.0725
R3051 VGND.n1110 VGND.n624 3.0725
R3052 VGND.n1111 VGND.n1110 3.0725
R3053 VGND.n1112 VGND.n1111 3.0725
R3054 VGND.n1112 VGND.n616 3.0725
R3055 VGND.n1122 VGND.n616 3.0725
R3056 VGND.n1123 VGND.n1122 3.0725
R3057 VGND.n1124 VGND.n1123 3.0725
R3058 VGND.n1124 VGND.n607 3.0725
R3059 VGND.n1134 VGND.n607 3.0725
R3060 VGND.n1135 VGND.n1134 3.0725
R3061 VGND.n1136 VGND.n1135 3.0725
R3062 VGND.n1136 VGND.n600 3.0725
R3063 VGND.n1146 VGND.n600 3.0725
R3064 VGND.n1147 VGND.n1146 3.0725
R3065 VGND.n1148 VGND.n1147 3.0725
R3066 VGND.n1148 VGND.n592 3.0725
R3067 VGND.n1158 VGND.n592 3.0725
R3068 VGND.n1159 VGND.n1158 3.0725
R3069 VGND.n1160 VGND.n1159 3.0725
R3070 VGND.n1160 VGND.n584 3.0725
R3071 VGND.n1170 VGND.n584 3.0725
R3072 VGND.n1171 VGND.n1170 3.0725
R3073 VGND.n1172 VGND.n1171 3.0725
R3074 VGND.n1172 VGND.n576 3.0725
R3075 VGND.n1182 VGND.n576 3.0725
R3076 VGND.n1183 VGND.n1182 3.0725
R3077 VGND.n1184 VGND.n1183 3.0725
R3078 VGND.n1184 VGND.n567 3.0725
R3079 VGND.n1194 VGND.n567 3.0725
R3080 VGND.n1195 VGND.n1194 3.0725
R3081 VGND.n1196 VGND.n1195 3.0725
R3082 VGND.n1196 VGND.n560 3.0725
R3083 VGND.n1206 VGND.n560 3.0725
R3084 VGND.n1207 VGND.n1206 3.0725
R3085 VGND.n1208 VGND.n1207 3.0725
R3086 VGND.n1208 VGND.n552 3.0725
R3087 VGND.n1218 VGND.n552 3.0725
R3088 VGND.n1219 VGND.n1218 3.0725
R3089 VGND.n1220 VGND.n1219 3.0725
R3090 VGND.n1220 VGND.n544 3.0725
R3091 VGND.n1230 VGND.n544 3.0725
R3092 VGND.n1231 VGND.n1230 3.0725
R3093 VGND.n1232 VGND.n1231 3.0725
R3094 VGND.n1232 VGND.n536 3.0725
R3095 VGND.n1242 VGND.n536 3.0725
R3096 VGND.n1243 VGND.n1242 3.0725
R3097 VGND.n1244 VGND.n1243 3.0725
R3098 VGND.n1244 VGND.n527 3.0725
R3099 VGND.n1254 VGND.n527 3.0725
R3100 VGND.n1255 VGND.n1254 3.0725
R3101 VGND.n1256 VGND.n1255 3.0725
R3102 VGND.n1256 VGND.n520 3.0725
R3103 VGND.n1266 VGND.n520 3.0725
R3104 VGND.n1267 VGND.n1266 3.0725
R3105 VGND.n1268 VGND.n1267 3.0725
R3106 VGND.n1268 VGND.n512 3.0725
R3107 VGND.n1278 VGND.n512 3.0725
R3108 VGND.n1279 VGND.n1278 3.0725
R3109 VGND.n1280 VGND.n1279 3.0725
R3110 VGND.n1280 VGND.n504 3.0725
R3111 VGND.n1290 VGND.n504 3.0725
R3112 VGND.n1291 VGND.n1290 3.0725
R3113 VGND.n1292 VGND.n1291 3.0725
R3114 VGND.n1292 VGND.n496 3.0725
R3115 VGND.n1302 VGND.n496 3.0725
R3116 VGND.n1303 VGND.n1302 3.0725
R3117 VGND.n1307 VGND.n1303 3.0725
R3118 VGND.n1307 VGND.n1306 3.0725
R3119 VGND.n1306 VGND.n1305 3.0725
R3120 VGND.n1305 VGND.n486 3.0725
R3121 VGND.n1476 VGND.n486 3.0725
R3122 VGND.n1476 VGND.n1475 3.0725
R3123 VGND.n1475 VGND.n1318 3.0725
R3124 VGND.n1471 VGND.n1318 3.0725
R3125 VGND.n1471 VGND.n1470 3.0725
R3126 VGND.n1470 VGND.n1469 3.0725
R3127 VGND.n1469 VGND.n1321 3.0725
R3128 VGND.n1465 VGND.n1321 3.0725
R3129 VGND.n1465 VGND.n1464 3.0725
R3130 VGND.n1464 VGND.n1463 3.0725
R3131 VGND.n1463 VGND.n1324 3.0725
R3132 VGND.n1459 VGND.n1324 3.0725
R3133 VGND.n1459 VGND.n1458 3.0725
R3134 VGND.n1458 VGND.n1457 3.0725
R3135 VGND.n1457 VGND.n1327 3.0725
R3136 VGND.n1453 VGND.n1327 3.0725
R3137 VGND.n1453 VGND.n1452 3.0725
R3138 VGND.n1452 VGND.n1451 3.0725
R3139 VGND.n1451 VGND.n1330 3.0725
R3140 VGND.n1447 VGND.n1330 3.0725
R3141 VGND.n1447 VGND.n1446 3.0725
R3142 VGND.n1446 VGND.n1445 3.0725
R3143 VGND.n1445 VGND.n1333 3.0725
R3144 VGND.n1441 VGND.n1333 3.0725
R3145 VGND.n1441 VGND.n1440 3.0725
R3146 VGND.n1440 VGND.n1439 3.0725
R3147 VGND.n1439 VGND.n1336 3.0725
R3148 VGND.n1435 VGND.n1336 3.0725
R3149 VGND.n1435 VGND.n1434 3.0725
R3150 VGND.n1434 VGND.n1433 3.0725
R3151 VGND.n1433 VGND.n1339 3.0725
R3152 VGND.n1429 VGND.n1339 3.0725
R3153 VGND.n1429 VGND.n1428 3.0725
R3154 VGND.n1428 VGND.n1427 3.0725
R3155 VGND.n1427 VGND.n1342 3.0725
R3156 VGND.n1423 VGND.n1342 3.0725
R3157 VGND.n1423 VGND.n1422 3.0725
R3158 VGND.n1422 VGND.n1421 3.0725
R3159 VGND.n1421 VGND.n1345 3.0725
R3160 VGND.n1417 VGND.n1345 3.0725
R3161 VGND.n1417 VGND.n1416 3.0725
R3162 VGND.n1416 VGND.n1415 3.0725
R3163 VGND.n1415 VGND.n1348 3.0725
R3164 VGND.n1411 VGND.n1348 3.0725
R3165 VGND.n1411 VGND.n1410 3.0725
R3166 VGND.n1410 VGND.n1409 3.0725
R3167 VGND.n1409 VGND.n1351 3.0725
R3168 VGND.n1405 VGND.n1351 3.0725
R3169 VGND.n1405 VGND.n1404 3.0725
R3170 VGND.n1404 VGND.n1403 3.0725
R3171 VGND.n1403 VGND.n1354 3.0725
R3172 VGND.n1399 VGND.n1354 3.0725
R3173 VGND.n1399 VGND.n1398 3.0725
R3174 VGND.n1398 VGND.n1397 3.0725
R3175 VGND.n1397 VGND.n1357 3.0725
R3176 VGND.n1393 VGND.n1357 3.0725
R3177 VGND.n1393 VGND.n1392 3.0725
R3178 VGND.n1392 VGND.n1391 3.0725
R3179 VGND.n1391 VGND.n1360 3.0725
R3180 VGND.n1387 VGND.n1360 3.0725
R3181 VGND.n1387 VGND.n1386 3.0725
R3182 VGND.n1386 VGND.n1385 3.0725
R3183 VGND.n1385 VGND.n1363 3.0725
R3184 VGND.n1381 VGND.n1363 3.0725
R3185 VGND.n1381 VGND.n1380 3.0725
R3186 VGND.n1380 VGND.n1379 3.0725
R3187 VGND.n1379 VGND.n1366 3.0725
R3188 VGND.n1375 VGND.n1366 3.0725
R3189 VGND.n1375 VGND.n1374 3.0725
R3190 VGND.n1374 VGND.n1373 3.0725
R3191 VGND.n1373 VGND.n1369 3.0725
R3192 VGND.n1369 VGND.n99 3.0725
R3193 VGND.n1563 VGND.n100 3.0725
R3194 VGND.n1559 VGND.n100 3.0725
R3195 VGND.n1559 VGND.n1558 3.0725
R3196 VGND.n1558 VGND.n1557 3.0725
R3197 VGND.n1557 VGND.n1556 3.0725
R3198 VGND.n1556 VGND.n1555 3.0725
R3199 VGND.n1555 VGND.n1554 3.0725
R3200 VGND.n1554 VGND.n1553 3.0725
R3201 VGND.n1553 VGND.n1552 3.0725
R3202 VGND.n1552 VGND.n1551 3.0725
R3203 VGND.n1551 VGND.n1550 3.0725
R3204 VGND.n1550 VGND.n1549 3.0725
R3205 VGND.n1549 VGND.n1548 3.0725
R3206 VGND.n1548 VGND.n1547 3.0725
R3207 VGND.n1547 VGND.n1546 3.0725
R3208 VGND.n1546 VGND.n1545 3.0725
R3209 VGND.n1545 VGND.n1544 3.0725
R3210 VGND.n1544 VGND.n1543 3.0725
R3211 VGND.n1543 VGND.n1542 3.0725
R3212 VGND.n1542 VGND.n1541 3.0725
R3213 VGND.n1541 VGND.n1540 3.0725
R3214 VGND.n1540 VGND.n1539 3.0725
R3215 VGND.n1539 VGND.n1538 3.0725
R3216 VGND.n1538 VGND.n1537 3.0725
R3217 VGND.n1537 VGND.n1536 3.0725
R3218 VGND.n1536 VGND.n1535 3.0725
R3219 VGND.n1535 VGND.n1534 3.0725
R3220 VGND.n1534 VGND.n1533 3.0725
R3221 VGND.n1533 VGND.n1532 3.0725
R3222 VGND.n1532 VGND.n1531 3.0725
R3223 VGND.n1531 VGND.n1530 3.0725
R3224 VGND.n1530 VGND.n1529 3.0725
R3225 VGND.n1529 VGND.n1528 3.0725
R3226 VGND.n1528 VGND.n1527 3.0725
R3227 VGND.n1527 VGND.n1526 3.0725
R3228 VGND.n1526 VGND.n1525 3.0725
R3229 VGND.n1525 VGND.n1524 3.0725
R3230 VGND.n1524 VGND.n1523 3.0725
R3231 VGND.n1523 VGND.n1522 3.0725
R3232 VGND.n1522 VGND.n1521 3.0725
R3233 VGND.n1521 VGND.n1520 3.0725
R3234 VGND.n1520 VGND.n1519 3.0725
R3235 VGND.n1519 VGND.n1518 3.0725
R3236 VGND.n1518 VGND.n1517 3.0725
R3237 VGND.n1517 VGND.n1516 3.0725
R3238 VGND.n1516 VGND.n1515 3.0725
R3239 VGND.n1515 VGND.n1514 3.0725
R3240 VGND.n1514 VGND.n1513 3.0725
R3241 VGND.n1513 VGND.n1512 3.0725
R3242 VGND.n1512 VGND.n1511 3.0725
R3243 VGND.n1511 VGND.n1510 3.0725
R3244 VGND.n1510 VGND.n1509 3.0725
R3245 VGND.n1509 VGND.n1508 3.0725
R3246 VGND.n1508 VGND.n1507 3.0725
R3247 VGND.n1507 VGND.n1506 3.0725
R3248 VGND.n1506 VGND.n1505 3.0725
R3249 VGND.n1505 VGND.n1504 3.0725
R3250 VGND.n1504 VGND.n1503 3.0725
R3251 VGND.n1503 VGND.n1502 3.0725
R3252 VGND.n1502 VGND.n1501 3.0725
R3253 VGND.n1501 VGND.n1500 3.0725
R3254 VGND.n1500 VGND.n1499 3.0725
R3255 VGND.n1499 VGND.n1498 3.0725
R3256 VGND.n1498 VGND.n1497 3.0725
R3257 VGND.n1497 VGND.n1496 3.0725
R3258 VGND.n1496 VGND.n1495 3.0725
R3259 VGND.n1495 VGND.n1494 3.0725
R3260 VGND.n1494 VGND.n1493 3.0725
R3261 VGND.n1493 VGND.n1492 3.0725
R3262 VGND.n1492 VGND.n1491 3.0725
R3263 VGND.n1491 VGND.n1490 3.0725
R3264 VGND.n1490 VGND.n1489 3.0725
R3265 VGND.n1489 VGND.n1488 3.0725
R3266 VGND.n1488 VGND.n1487 3.0725
R3267 VGND.n1487 VGND.n1486 3.0725
R3268 VGND.n1486 VGND.n1485 3.0725
R3269 VGND.n484 VGND.n483 3.0725
R3270 VGND.n483 VGND.n482 3.0725
R3271 VGND.n482 VGND.n481 3.0725
R3272 VGND.n481 VGND.n480 3.0725
R3273 VGND.n480 VGND.n479 3.0725
R3274 VGND.n479 VGND.n478 3.0725
R3275 VGND.n478 VGND.n477 3.0725
R3276 VGND.n477 VGND.n476 3.0725
R3277 VGND.n476 VGND.n475 3.0725
R3278 VGND.n475 VGND.n474 3.0725
R3279 VGND.n474 VGND.n473 3.0725
R3280 VGND.n473 VGND.n472 3.0725
R3281 VGND.n472 VGND.n471 3.0725
R3282 VGND.n471 VGND.n470 3.0725
R3283 VGND.n470 VGND.n469 3.0725
R3284 VGND.n469 VGND.n468 3.0725
R3285 VGND.n468 VGND.n467 3.0725
R3286 VGND.n467 VGND.n466 3.0725
R3287 VGND.n466 VGND.n465 3.0725
R3288 VGND.n465 VGND.n464 3.0725
R3289 VGND.n464 VGND.n463 3.0725
R3290 VGND.n463 VGND.n462 3.0725
R3291 VGND.n462 VGND.n461 3.0725
R3292 VGND.n461 VGND.n460 3.0725
R3293 VGND.n460 VGND.n459 3.0725
R3294 VGND.n459 VGND.n458 3.0725
R3295 VGND.n458 VGND.n457 3.0725
R3296 VGND.n457 VGND.n456 3.0725
R3297 VGND.n456 VGND.n455 3.0725
R3298 VGND.n455 VGND.n454 3.0725
R3299 VGND.n454 VGND.n453 3.0725
R3300 VGND.n453 VGND.n452 3.0725
R3301 VGND.n452 VGND.n451 3.0725
R3302 VGND.n451 VGND.n450 3.0725
R3303 VGND.n450 VGND.n449 3.0725
R3304 VGND.n449 VGND.n448 3.0725
R3305 VGND.n448 VGND.n447 3.0725
R3306 VGND.n447 VGND.n446 3.0725
R3307 VGND.n446 VGND.n445 3.0725
R3308 VGND.n445 VGND.n444 3.0725
R3309 VGND.n444 VGND.n443 3.0725
R3310 VGND.n443 VGND.n442 3.0725
R3311 VGND.n442 VGND.n441 3.0725
R3312 VGND.n441 VGND.n440 3.0725
R3313 VGND.n440 VGND.n439 3.0725
R3314 VGND.n439 VGND.n438 3.0725
R3315 VGND.n438 VGND.n437 3.0725
R3316 VGND.n437 VGND.n436 3.0725
R3317 VGND.n436 VGND.n435 3.0725
R3318 VGND.n435 VGND.n434 3.0725
R3319 VGND.n434 VGND.n433 3.0725
R3320 VGND.n433 VGND.n432 3.0725
R3321 VGND.n432 VGND.n431 3.0725
R3322 VGND.n431 VGND.n430 3.0725
R3323 VGND.n430 VGND.n429 3.0725
R3324 VGND.n429 VGND.n428 3.0725
R3325 VGND.n428 VGND.n427 3.0725
R3326 VGND.n427 VGND.n426 3.0725
R3327 VGND.n426 VGND.n425 3.0725
R3328 VGND.n425 VGND.n424 3.0725
R3329 VGND.n424 VGND.n423 3.0725
R3330 VGND.n423 VGND.n422 3.0725
R3331 VGND.n422 VGND.n421 3.0725
R3332 VGND.n421 VGND.n420 3.0725
R3333 VGND.n420 VGND.n419 3.0725
R3334 VGND.n419 VGND.n418 3.0725
R3335 VGND.n418 VGND.n417 3.0725
R3336 VGND.n417 VGND.n416 3.0725
R3337 VGND.n416 VGND.n415 3.0725
R3338 VGND.n415 VGND.n414 3.0725
R3339 VGND.n414 VGND.n413 3.0725
R3340 VGND.n413 VGND.n412 3.0725
R3341 VGND.n412 VGND.n411 3.0725
R3342 VGND.n411 VGND.n410 3.0725
R3343 VGND.n410 VGND.n409 3.0725
R3344 VGND.n409 VGND.n94 3.0725
R3345 VGND.n1106 VGND.n1105 3.0725
R3346 VGND.n1106 VGND.n620 3.0725
R3347 VGND.n1116 VGND.n620 3.0725
R3348 VGND.n1117 VGND.n1116 3.0725
R3349 VGND.n1118 VGND.n1117 3.0725
R3350 VGND.n1118 VGND.n612 3.0725
R3351 VGND.n1128 VGND.n612 3.0725
R3352 VGND.n1129 VGND.n1128 3.0725
R3353 VGND.n1130 VGND.n1129 3.0725
R3354 VGND.n1130 VGND.n604 3.0725
R3355 VGND.n1140 VGND.n604 3.0725
R3356 VGND.n1141 VGND.n1140 3.0725
R3357 VGND.n1142 VGND.n1141 3.0725
R3358 VGND.n1142 VGND.n596 3.0725
R3359 VGND.n1152 VGND.n596 3.0725
R3360 VGND.n1153 VGND.n1152 3.0725
R3361 VGND.n1154 VGND.n1153 3.0725
R3362 VGND.n1154 VGND.n587 3.0725
R3363 VGND.n1164 VGND.n587 3.0725
R3364 VGND.n1165 VGND.n1164 3.0725
R3365 VGND.n1166 VGND.n1165 3.0725
R3366 VGND.n1166 VGND.n580 3.0725
R3367 VGND.n1176 VGND.n580 3.0725
R3368 VGND.n1177 VGND.n1176 3.0725
R3369 VGND.n1178 VGND.n1177 3.0725
R3370 VGND.n1178 VGND.n572 3.0725
R3371 VGND.n1188 VGND.n572 3.0725
R3372 VGND.n1189 VGND.n1188 3.0725
R3373 VGND.n1190 VGND.n1189 3.0725
R3374 VGND.n1190 VGND.n564 3.0725
R3375 VGND.n1200 VGND.n564 3.0725
R3376 VGND.n1201 VGND.n1200 3.0725
R3377 VGND.n1202 VGND.n1201 3.0725
R3378 VGND.n1202 VGND.n556 3.0725
R3379 VGND.n1212 VGND.n556 3.0725
R3380 VGND.n1213 VGND.n1212 3.0725
R3381 VGND.n1214 VGND.n1213 3.0725
R3382 VGND.n1214 VGND.n547 3.0725
R3383 VGND.n1224 VGND.n547 3.0725
R3384 VGND.n1225 VGND.n1224 3.0725
R3385 VGND.n1226 VGND.n1225 3.0725
R3386 VGND.n1226 VGND.n540 3.0725
R3387 VGND.n1236 VGND.n540 3.0725
R3388 VGND.n1237 VGND.n1236 3.0725
R3389 VGND.n1238 VGND.n1237 3.0725
R3390 VGND.n1238 VGND.n532 3.0725
R3391 VGND.n1248 VGND.n532 3.0725
R3392 VGND.n1249 VGND.n1248 3.0725
R3393 VGND.n1250 VGND.n1249 3.0725
R3394 VGND.n1250 VGND.n524 3.0725
R3395 VGND.n1260 VGND.n524 3.0725
R3396 VGND.n1261 VGND.n1260 3.0725
R3397 VGND.n1262 VGND.n1261 3.0725
R3398 VGND.n1262 VGND.n516 3.0725
R3399 VGND.n1272 VGND.n516 3.0725
R3400 VGND.n1273 VGND.n1272 3.0725
R3401 VGND.n1274 VGND.n1273 3.0725
R3402 VGND.n1274 VGND.n507 3.0725
R3403 VGND.n1284 VGND.n507 3.0725
R3404 VGND.n1285 VGND.n1284 3.0725
R3405 VGND.n1286 VGND.n1285 3.0725
R3406 VGND.n1286 VGND.n500 3.0725
R3407 VGND.n1296 VGND.n500 3.0725
R3408 VGND.n1297 VGND.n1296 3.0725
R3409 VGND.n1298 VGND.n1297 3.0725
R3410 VGND.n1298 VGND.n490 3.0725
R3411 VGND.n1311 VGND.n490 3.0725
R3412 VGND.n1312 VGND.n1311 3.0725
R3413 VGND.n1313 VGND.n1312 3.0725
R3414 VGND.n1313 VGND.n2 3.0725
R3415 VGND.n1676 VGND.n2 3.0725
R3416 VGND.n1676 VGND.n1675 3.0725
R3417 VGND.n1675 VGND.n4 3.0725
R3418 VGND.n1671 VGND.n4 3.0725
R3419 VGND.n1671 VGND.n1670 3.0725
R3420 VGND.n1670 VGND.n1669 3.0725
R3421 VGND.n1669 VGND.n9 3.0725
R3422 VGND.n1665 VGND.n9 3.0725
R3423 VGND.n1665 VGND.n1664 3.0725
R3424 VGND.n1664 VGND.n1663 3.0725
R3425 VGND.n1663 VGND.n14 3.0725
R3426 VGND.n1659 VGND.n14 3.0725
R3427 VGND.n1659 VGND.n1658 3.0725
R3428 VGND.n1658 VGND.n1657 3.0725
R3429 VGND.n1657 VGND.n19 3.0725
R3430 VGND.n1653 VGND.n19 3.0725
R3431 VGND.n1653 VGND.n1652 3.0725
R3432 VGND.n1652 VGND.n1651 3.0725
R3433 VGND.n1651 VGND.n24 3.0725
R3434 VGND.n1647 VGND.n24 3.0725
R3435 VGND.n1647 VGND.n1646 3.0725
R3436 VGND.n1646 VGND.n1645 3.0725
R3437 VGND.n1645 VGND.n29 3.0725
R3438 VGND.n1641 VGND.n29 3.0725
R3439 VGND.n1641 VGND.n1640 3.0725
R3440 VGND.n1640 VGND.n1639 3.0725
R3441 VGND.n1639 VGND.n34 3.0725
R3442 VGND.n1635 VGND.n34 3.0725
R3443 VGND.n1635 VGND.n1634 3.0725
R3444 VGND.n1634 VGND.n1633 3.0725
R3445 VGND.n1633 VGND.n39 3.0725
R3446 VGND.n1629 VGND.n39 3.0725
R3447 VGND.n1629 VGND.n1628 3.0725
R3448 VGND.n1628 VGND.n1627 3.0725
R3449 VGND.n1627 VGND.n44 3.0725
R3450 VGND.n1623 VGND.n44 3.0725
R3451 VGND.n1623 VGND.n1622 3.0725
R3452 VGND.n1622 VGND.n1621 3.0725
R3453 VGND.n1621 VGND.n49 3.0725
R3454 VGND.n1617 VGND.n49 3.0725
R3455 VGND.n1617 VGND.n1616 3.0725
R3456 VGND.n1616 VGND.n1615 3.0725
R3457 VGND.n1615 VGND.n54 3.0725
R3458 VGND.n1611 VGND.n54 3.0725
R3459 VGND.n1611 VGND.n1610 3.0725
R3460 VGND.n1610 VGND.n1609 3.0725
R3461 VGND.n1609 VGND.n59 3.0725
R3462 VGND.n1605 VGND.n59 3.0725
R3463 VGND.n1605 VGND.n1604 3.0725
R3464 VGND.n1604 VGND.n1603 3.0725
R3465 VGND.n1603 VGND.n64 3.0725
R3466 VGND.n1599 VGND.n64 3.0725
R3467 VGND.n1599 VGND.n1598 3.0725
R3468 VGND.n1598 VGND.n1597 3.0725
R3469 VGND.n1597 VGND.n69 3.0725
R3470 VGND.n1593 VGND.n69 3.0725
R3471 VGND.n1593 VGND.n1592 3.0725
R3472 VGND.n1592 VGND.n1591 3.0725
R3473 VGND.n1591 VGND.n74 3.0725
R3474 VGND.n1587 VGND.n74 3.0725
R3475 VGND.n1587 VGND.n1586 3.0725
R3476 VGND.n1586 VGND.n1585 3.0725
R3477 VGND.n1585 VGND.n79 3.0725
R3478 VGND.n1581 VGND.n79 3.0725
R3479 VGND.n1581 VGND.n1580 3.0725
R3480 VGND.n1580 VGND.n1579 3.0725
R3481 VGND.n1579 VGND.n84 3.0725
R3482 VGND.n1575 VGND.n84 3.0725
R3483 VGND.n1575 VGND.n1574 3.0725
R3484 VGND.n1574 VGND.n1573 3.0725
R3485 VGND.n1573 VGND.n89 3.0725
R3486 VGND.n1569 VGND.n89 3.0725
R3487 VGND.n1258 VGND.t13 2.97046
R3488 VGND.n1331 VGND.t7 2.97046
R3489 VGND.t26 VGND.n514 2.22797
R3490 VGND.t16 VGND.n22 2.22797
R3491 VGND.n1677 VGND.n1 2.21883
R3492 VGND.n1477 VGND.n485 2.21883
R3493 VGND VGND.n1677 2.14633
R3494 VGND.n1019 VGND.n485 2.08592
R3495 VGND.n1019 VGND.n1 2.08592
R3496 VGND.n1483 VGND.n1481 2.08592
R3497 VGND.n1483 VGND.n1482 2.08592
R3498 VGND.n1481 VGND 1.82895
R3499 VGND.n942 VGND.n624 1.62183
R3500 VGND.n1564 VGND.n99 1.62183
R3501 VGND.n1105 VGND.n1104 1.62183
R3502 VGND.n1569 VGND.n1568 1.62183
R3503 VGND.n1021 VGND.n1020 1.5365
R3504 VGND.n1020 VGND.n1018 1.5365
R3505 VGND.n1485 VGND.n1484 1.5365
R3506 VGND.n1484 VGND.n484 1.5365
R3507 VGND.n1288 VGND.t1 1.48548
R3508 VGND.t29 VGND.n16 1.48548
R3509 VGND.n1478 VGND.n1477 1.358
R3510 VGND.n1478 VGND.t18 0.952889
R3511 VGND.n485 VGND.t9 0.901512
R3512 VGND.n1 VGND.t10 0.901501
R3513 VGND.n1479 VGND.n1478 0.861333
R3514 VGND.n1480 VGND.t24 0.769683
R3515 VGND.n0 VGND.t25 0.769672
R3516 VGND.n1099 VGND.n629 0.742991
R3517 VGND.n632 VGND.n630 0.742991
R3518 VGND.n938 VGND.n937 0.742991
R3519 VGND.n1108 VGND.n626 0.742991
R3520 VGND.t22 VGND.n492 0.742991
R3521 VGND.t27 VGND.n10 0.742991
R3522 VGND.n103 VGND.n91 0.742991
R3523 VGND.n1561 VGND.n92 0.742991
R3524 VGND.n181 VGND.n96 0.742991
R3525 VGND.n1566 VGND.n97 0.742991
R3526 VGND.n1482 VGND 0.248417
R3527 VGND.n1678 VGND 0.073
R3528 VGND.n1481 VGND.n1480 0.0368793
R3529 VGND.n1678 VGND.n0 0.0368793
R3530 VGND.n1480 VGND.n1479 0.0367069
R3531 VGND.n1482 VGND.n0 0.0367069
R3532 VGND VGND.n1678 0.0305
R3533 VGND.n1677 VGND.n1676 0.0163163
R3534 VGND.n1477 VGND.n1476 0.0163163
R3535 VGND.n1020 VGND.n1019 0.0155974
R3536 VGND.n1484 VGND.n1483 0.0155974
R3537 D1 D1.t0 1.05785
R3538 OUT.n0 OUT.t0 0.823424
R3539 OUT.n0 OUT.t1 0.823424
R3540 OUT OUT.n0 0.17647
R3541 D2 D2.t0 1.05785
R3542 D3 D3.t0 1.05785
R3543 D4 D4.t0 1.05785
R3544 D5 D5.t0 1.05785
R3545 D6 D6.t0 1.05785
R3546 D0 D0.t0 1.05785
R3547 D7 D7.t0 1.05785
C0 a_840_493# a_1564_493# 0.337752f
C1 a_5908_493# a_4460_10921# 0.338797f
C2 D2 a_3374_10921# 0.389424f
C3 D1 a_3374_10921# 0.388627f
C4 D4 D3 0.024257f
C5 a_5546_10921# D3 0.388627f
C6 D2 a_4460_10921# 0.388627f
C7 a_9166_493# a_7718_10921# 0.338797f
C8 a_1202_10921# a_1564_493# 0.338797f
C9 D0 a_1202_10921# 0.388627f
C10 D3 a_4460_10921# 0.389424f
C11 a_2288_10921# a_3374_10921# 0.569962f
C12 a_6632_10921# a_7718_10921# 0.569962f
C13 a_3736_493# a_3374_10921# 0.338797f
C14 D1 D2 0.024257f
C15 a_6994_493# a_6632_10921# 0.338797f
C16 a_2650_493# a_1202_10921# 0.338797f
C17 OUT D7 0.473447f
C18 D2 D3 0.024257f
C19 D6 D5 0.024257f
C20 a_8080_493# a_7718_10921# 0.338797f
C21 a_6994_493# a_5546_10921# 0.338797f
C22 a_4822_493# a_3374_10921# 0.338797f
C23 a_2650_493# a_2288_10921# 0.338797f
C24 a_2288_10921# D1 0.389424f
C25 a_2288_10921# a_1202_10921# 0.569962f
C26 D4 a_6632_10921# 0.388627f
C27 D5 a_7718_10921# 0.388627f
C28 a_6632_10921# a_5546_10921# 0.569962f
C29 a_4822_493# a_4460_10921# 0.338797f
C30 a_8080_493# a_6632_10921# 0.338797f
C31 D4 a_5546_10921# 0.389424f
C32 D5 a_6632_10921# 0.389424f
C33 a_2288_10921# a_3736_493# 0.338797f
C34 D6 OUT 0.473447f
C35 a_5546_10921# a_4460_10921# 0.569962f
C36 a_3374_10921# a_4460_10921# 0.569962f
C37 a_5546_10921# a_5908_493# 0.338797f
C38 D4 D5 0.024257f
C39 D6 a_7718_10921# 0.389424f
C40 D7 VGND 0.882964f
C41 OUT VGND 0.991791f
C42 D6 VGND 0.465536f
C43 D5 VGND 0.46853f
C44 D4 VGND 0.46853f
C45 D3 VGND 0.46853f
C46 D2 VGND 0.46853f
C47 D1 VGND 0.489659f
C48 D0 VGND 0.906593f
C49 a_9166_493# VGND 1.18199f
C50 a_8080_493# VGND 0.844742f
C51 a_7718_10921# VGND 4.89913f
C52 a_6994_493# VGND 0.845481f
C53 a_6632_10921# VGND 4.31982f
C54 a_5908_493# VGND 0.845481f
C55 a_5546_10921# VGND 4.31982f
C56 a_4822_493# VGND 0.845481f
C57 a_4460_10921# VGND 4.31982f
C58 a_3736_493# VGND 0.845481f
C59 a_3374_10921# VGND 4.319839f
C60 a_2650_493# VGND 0.845481f
C61 a_2288_10921# VGND 4.65815f
C62 a_1564_493# VGND 0.844286f
C63 a_1202_10921# VGND 5.23785f
C64 a_840_493# VGND 1.18199f
.ends

